magic
tech sky130A
magscale 1 2
timestamp 1652625669
<< obsli1 >>
rect 1104 2159 148856 47345
<< obsm1 >>
rect 106 1844 149762 47376
<< metal2 >>
rect 2778 49200 2834 50000
rect 8298 49200 8354 50000
rect 13818 49200 13874 50000
rect 19430 49200 19486 50000
rect 24950 49200 25006 50000
rect 30470 49200 30526 50000
rect 36082 49200 36138 50000
rect 41602 49200 41658 50000
rect 47122 49200 47178 50000
rect 52734 49200 52790 50000
rect 58254 49200 58310 50000
rect 63866 49200 63922 50000
rect 69386 49200 69442 50000
rect 74906 49200 74962 50000
rect 80518 49200 80574 50000
rect 86038 49200 86094 50000
rect 91558 49200 91614 50000
rect 97170 49200 97226 50000
rect 102690 49200 102746 50000
rect 108302 49200 108358 50000
rect 113822 49200 113878 50000
rect 119342 49200 119398 50000
rect 124954 49200 125010 50000
rect 130474 49200 130530 50000
rect 135994 49200 136050 50000
rect 141606 49200 141662 50000
rect 147126 49200 147182 50000
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123850 0 123906 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124770 0 124826 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130290 0 130346 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131762 0 131818 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135442 0 135498 800
rect 135718 0 135774 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138478 0 138534 800
rect 138754 0 138810 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142434 0 142490 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143630 0 143686 800
rect 143906 0 143962 800
rect 144274 0 144330 800
rect 144550 0 144606 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146666 0 146722 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147586 0 147642 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149426 0 149482 800
rect 149702 0 149758 800
<< obsm2 >>
rect 112 49144 2722 49473
rect 2890 49144 8242 49473
rect 8410 49144 13762 49473
rect 13930 49144 19374 49473
rect 19542 49144 24894 49473
rect 25062 49144 30414 49473
rect 30582 49144 36026 49473
rect 36194 49144 41546 49473
rect 41714 49144 47066 49473
rect 47234 49144 52678 49473
rect 52846 49144 58198 49473
rect 58366 49144 63810 49473
rect 63978 49144 69330 49473
rect 69498 49144 74850 49473
rect 75018 49144 80462 49473
rect 80630 49144 85982 49473
rect 86150 49144 91502 49473
rect 91670 49144 97114 49473
rect 97282 49144 102634 49473
rect 102802 49144 108246 49473
rect 108414 49144 113766 49473
rect 113934 49144 119286 49473
rect 119454 49144 124898 49473
rect 125066 49144 130418 49473
rect 130586 49144 135938 49473
rect 136106 49144 141550 49473
rect 141718 49144 147070 49473
rect 147238 49144 149756 49473
rect 112 856 149756 49144
rect 222 575 330 856
rect 498 575 606 856
rect 774 575 882 856
rect 1050 575 1250 856
rect 1418 575 1526 856
rect 1694 575 1802 856
rect 1970 575 2170 856
rect 2338 575 2446 856
rect 2614 575 2722 856
rect 2890 575 3090 856
rect 3258 575 3366 856
rect 3534 575 3642 856
rect 3810 575 3918 856
rect 4086 575 4286 856
rect 4454 575 4562 856
rect 4730 575 4838 856
rect 5006 575 5206 856
rect 5374 575 5482 856
rect 5650 575 5758 856
rect 5926 575 6126 856
rect 6294 575 6402 856
rect 6570 575 6678 856
rect 6846 575 7046 856
rect 7214 575 7322 856
rect 7490 575 7598 856
rect 7766 575 7874 856
rect 8042 575 8242 856
rect 8410 575 8518 856
rect 8686 575 8794 856
rect 8962 575 9162 856
rect 9330 575 9438 856
rect 9606 575 9714 856
rect 9882 575 10082 856
rect 10250 575 10358 856
rect 10526 575 10634 856
rect 10802 575 11002 856
rect 11170 575 11278 856
rect 11446 575 11554 856
rect 11722 575 11830 856
rect 11998 575 12198 856
rect 12366 575 12474 856
rect 12642 575 12750 856
rect 12918 575 13118 856
rect 13286 575 13394 856
rect 13562 575 13670 856
rect 13838 575 14038 856
rect 14206 575 14314 856
rect 14482 575 14590 856
rect 14758 575 14958 856
rect 15126 575 15234 856
rect 15402 575 15510 856
rect 15678 575 15786 856
rect 15954 575 16154 856
rect 16322 575 16430 856
rect 16598 575 16706 856
rect 16874 575 17074 856
rect 17242 575 17350 856
rect 17518 575 17626 856
rect 17794 575 17994 856
rect 18162 575 18270 856
rect 18438 575 18546 856
rect 18714 575 18822 856
rect 18990 575 19190 856
rect 19358 575 19466 856
rect 19634 575 19742 856
rect 19910 575 20110 856
rect 20278 575 20386 856
rect 20554 575 20662 856
rect 20830 575 21030 856
rect 21198 575 21306 856
rect 21474 575 21582 856
rect 21750 575 21950 856
rect 22118 575 22226 856
rect 22394 575 22502 856
rect 22670 575 22778 856
rect 22946 575 23146 856
rect 23314 575 23422 856
rect 23590 575 23698 856
rect 23866 575 24066 856
rect 24234 575 24342 856
rect 24510 575 24618 856
rect 24786 575 24986 856
rect 25154 575 25262 856
rect 25430 575 25538 856
rect 25706 575 25906 856
rect 26074 575 26182 856
rect 26350 575 26458 856
rect 26626 575 26734 856
rect 26902 575 27102 856
rect 27270 575 27378 856
rect 27546 575 27654 856
rect 27822 575 28022 856
rect 28190 575 28298 856
rect 28466 575 28574 856
rect 28742 575 28942 856
rect 29110 575 29218 856
rect 29386 575 29494 856
rect 29662 575 29862 856
rect 30030 575 30138 856
rect 30306 575 30414 856
rect 30582 575 30690 856
rect 30858 575 31058 856
rect 31226 575 31334 856
rect 31502 575 31610 856
rect 31778 575 31978 856
rect 32146 575 32254 856
rect 32422 575 32530 856
rect 32698 575 32898 856
rect 33066 575 33174 856
rect 33342 575 33450 856
rect 33618 575 33726 856
rect 33894 575 34094 856
rect 34262 575 34370 856
rect 34538 575 34646 856
rect 34814 575 35014 856
rect 35182 575 35290 856
rect 35458 575 35566 856
rect 35734 575 35934 856
rect 36102 575 36210 856
rect 36378 575 36486 856
rect 36654 575 36854 856
rect 37022 575 37130 856
rect 37298 575 37406 856
rect 37574 575 37682 856
rect 37850 575 38050 856
rect 38218 575 38326 856
rect 38494 575 38602 856
rect 38770 575 38970 856
rect 39138 575 39246 856
rect 39414 575 39522 856
rect 39690 575 39890 856
rect 40058 575 40166 856
rect 40334 575 40442 856
rect 40610 575 40810 856
rect 40978 575 41086 856
rect 41254 575 41362 856
rect 41530 575 41638 856
rect 41806 575 42006 856
rect 42174 575 42282 856
rect 42450 575 42558 856
rect 42726 575 42926 856
rect 43094 575 43202 856
rect 43370 575 43478 856
rect 43646 575 43846 856
rect 44014 575 44122 856
rect 44290 575 44398 856
rect 44566 575 44766 856
rect 44934 575 45042 856
rect 45210 575 45318 856
rect 45486 575 45594 856
rect 45762 575 45962 856
rect 46130 575 46238 856
rect 46406 575 46514 856
rect 46682 575 46882 856
rect 47050 575 47158 856
rect 47326 575 47434 856
rect 47602 575 47802 856
rect 47970 575 48078 856
rect 48246 575 48354 856
rect 48522 575 48722 856
rect 48890 575 48998 856
rect 49166 575 49274 856
rect 49442 575 49550 856
rect 49718 575 49918 856
rect 50086 575 50194 856
rect 50362 575 50470 856
rect 50638 575 50838 856
rect 51006 575 51114 856
rect 51282 575 51390 856
rect 51558 575 51758 856
rect 51926 575 52034 856
rect 52202 575 52310 856
rect 52478 575 52586 856
rect 52754 575 52954 856
rect 53122 575 53230 856
rect 53398 575 53506 856
rect 53674 575 53874 856
rect 54042 575 54150 856
rect 54318 575 54426 856
rect 54594 575 54794 856
rect 54962 575 55070 856
rect 55238 575 55346 856
rect 55514 575 55714 856
rect 55882 575 55990 856
rect 56158 575 56266 856
rect 56434 575 56542 856
rect 56710 575 56910 856
rect 57078 575 57186 856
rect 57354 575 57462 856
rect 57630 575 57830 856
rect 57998 575 58106 856
rect 58274 575 58382 856
rect 58550 575 58750 856
rect 58918 575 59026 856
rect 59194 575 59302 856
rect 59470 575 59670 856
rect 59838 575 59946 856
rect 60114 575 60222 856
rect 60390 575 60498 856
rect 60666 575 60866 856
rect 61034 575 61142 856
rect 61310 575 61418 856
rect 61586 575 61786 856
rect 61954 575 62062 856
rect 62230 575 62338 856
rect 62506 575 62706 856
rect 62874 575 62982 856
rect 63150 575 63258 856
rect 63426 575 63626 856
rect 63794 575 63902 856
rect 64070 575 64178 856
rect 64346 575 64454 856
rect 64622 575 64822 856
rect 64990 575 65098 856
rect 65266 575 65374 856
rect 65542 575 65742 856
rect 65910 575 66018 856
rect 66186 575 66294 856
rect 66462 575 66662 856
rect 66830 575 66938 856
rect 67106 575 67214 856
rect 67382 575 67490 856
rect 67658 575 67858 856
rect 68026 575 68134 856
rect 68302 575 68410 856
rect 68578 575 68778 856
rect 68946 575 69054 856
rect 69222 575 69330 856
rect 69498 575 69698 856
rect 69866 575 69974 856
rect 70142 575 70250 856
rect 70418 575 70618 856
rect 70786 575 70894 856
rect 71062 575 71170 856
rect 71338 575 71446 856
rect 71614 575 71814 856
rect 71982 575 72090 856
rect 72258 575 72366 856
rect 72534 575 72734 856
rect 72902 575 73010 856
rect 73178 575 73286 856
rect 73454 575 73654 856
rect 73822 575 73930 856
rect 74098 575 74206 856
rect 74374 575 74574 856
rect 74742 575 74850 856
rect 75018 575 75126 856
rect 75294 575 75402 856
rect 75570 575 75770 856
rect 75938 575 76046 856
rect 76214 575 76322 856
rect 76490 575 76690 856
rect 76858 575 76966 856
rect 77134 575 77242 856
rect 77410 575 77610 856
rect 77778 575 77886 856
rect 78054 575 78162 856
rect 78330 575 78530 856
rect 78698 575 78806 856
rect 78974 575 79082 856
rect 79250 575 79358 856
rect 79526 575 79726 856
rect 79894 575 80002 856
rect 80170 575 80278 856
rect 80446 575 80646 856
rect 80814 575 80922 856
rect 81090 575 81198 856
rect 81366 575 81566 856
rect 81734 575 81842 856
rect 82010 575 82118 856
rect 82286 575 82486 856
rect 82654 575 82762 856
rect 82930 575 83038 856
rect 83206 575 83314 856
rect 83482 575 83682 856
rect 83850 575 83958 856
rect 84126 575 84234 856
rect 84402 575 84602 856
rect 84770 575 84878 856
rect 85046 575 85154 856
rect 85322 575 85522 856
rect 85690 575 85798 856
rect 85966 575 86074 856
rect 86242 575 86350 856
rect 86518 575 86718 856
rect 86886 575 86994 856
rect 87162 575 87270 856
rect 87438 575 87638 856
rect 87806 575 87914 856
rect 88082 575 88190 856
rect 88358 575 88558 856
rect 88726 575 88834 856
rect 89002 575 89110 856
rect 89278 575 89478 856
rect 89646 575 89754 856
rect 89922 575 90030 856
rect 90198 575 90306 856
rect 90474 575 90674 856
rect 90842 575 90950 856
rect 91118 575 91226 856
rect 91394 575 91594 856
rect 91762 575 91870 856
rect 92038 575 92146 856
rect 92314 575 92514 856
rect 92682 575 92790 856
rect 92958 575 93066 856
rect 93234 575 93434 856
rect 93602 575 93710 856
rect 93878 575 93986 856
rect 94154 575 94262 856
rect 94430 575 94630 856
rect 94798 575 94906 856
rect 95074 575 95182 856
rect 95350 575 95550 856
rect 95718 575 95826 856
rect 95994 575 96102 856
rect 96270 575 96470 856
rect 96638 575 96746 856
rect 96914 575 97022 856
rect 97190 575 97390 856
rect 97558 575 97666 856
rect 97834 575 97942 856
rect 98110 575 98218 856
rect 98386 575 98586 856
rect 98754 575 98862 856
rect 99030 575 99138 856
rect 99306 575 99506 856
rect 99674 575 99782 856
rect 99950 575 100058 856
rect 100226 575 100426 856
rect 100594 575 100702 856
rect 100870 575 100978 856
rect 101146 575 101254 856
rect 101422 575 101622 856
rect 101790 575 101898 856
rect 102066 575 102174 856
rect 102342 575 102542 856
rect 102710 575 102818 856
rect 102986 575 103094 856
rect 103262 575 103462 856
rect 103630 575 103738 856
rect 103906 575 104014 856
rect 104182 575 104382 856
rect 104550 575 104658 856
rect 104826 575 104934 856
rect 105102 575 105210 856
rect 105378 575 105578 856
rect 105746 575 105854 856
rect 106022 575 106130 856
rect 106298 575 106498 856
rect 106666 575 106774 856
rect 106942 575 107050 856
rect 107218 575 107418 856
rect 107586 575 107694 856
rect 107862 575 107970 856
rect 108138 575 108338 856
rect 108506 575 108614 856
rect 108782 575 108890 856
rect 109058 575 109166 856
rect 109334 575 109534 856
rect 109702 575 109810 856
rect 109978 575 110086 856
rect 110254 575 110454 856
rect 110622 575 110730 856
rect 110898 575 111006 856
rect 111174 575 111374 856
rect 111542 575 111650 856
rect 111818 575 111926 856
rect 112094 575 112294 856
rect 112462 575 112570 856
rect 112738 575 112846 856
rect 113014 575 113122 856
rect 113290 575 113490 856
rect 113658 575 113766 856
rect 113934 575 114042 856
rect 114210 575 114410 856
rect 114578 575 114686 856
rect 114854 575 114962 856
rect 115130 575 115330 856
rect 115498 575 115606 856
rect 115774 575 115882 856
rect 116050 575 116250 856
rect 116418 575 116526 856
rect 116694 575 116802 856
rect 116970 575 117078 856
rect 117246 575 117446 856
rect 117614 575 117722 856
rect 117890 575 117998 856
rect 118166 575 118366 856
rect 118534 575 118642 856
rect 118810 575 118918 856
rect 119086 575 119286 856
rect 119454 575 119562 856
rect 119730 575 119838 856
rect 120006 575 120114 856
rect 120282 575 120482 856
rect 120650 575 120758 856
rect 120926 575 121034 856
rect 121202 575 121402 856
rect 121570 575 121678 856
rect 121846 575 121954 856
rect 122122 575 122322 856
rect 122490 575 122598 856
rect 122766 575 122874 856
rect 123042 575 123242 856
rect 123410 575 123518 856
rect 123686 575 123794 856
rect 123962 575 124070 856
rect 124238 575 124438 856
rect 124606 575 124714 856
rect 124882 575 124990 856
rect 125158 575 125358 856
rect 125526 575 125634 856
rect 125802 575 125910 856
rect 126078 575 126278 856
rect 126446 575 126554 856
rect 126722 575 126830 856
rect 126998 575 127198 856
rect 127366 575 127474 856
rect 127642 575 127750 856
rect 127918 575 128026 856
rect 128194 575 128394 856
rect 128562 575 128670 856
rect 128838 575 128946 856
rect 129114 575 129314 856
rect 129482 575 129590 856
rect 129758 575 129866 856
rect 130034 575 130234 856
rect 130402 575 130510 856
rect 130678 575 130786 856
rect 130954 575 131154 856
rect 131322 575 131430 856
rect 131598 575 131706 856
rect 131874 575 131982 856
rect 132150 575 132350 856
rect 132518 575 132626 856
rect 132794 575 132902 856
rect 133070 575 133270 856
rect 133438 575 133546 856
rect 133714 575 133822 856
rect 133990 575 134190 856
rect 134358 575 134466 856
rect 134634 575 134742 856
rect 134910 575 135018 856
rect 135186 575 135386 856
rect 135554 575 135662 856
rect 135830 575 135938 856
rect 136106 575 136306 856
rect 136474 575 136582 856
rect 136750 575 136858 856
rect 137026 575 137226 856
rect 137394 575 137502 856
rect 137670 575 137778 856
rect 137946 575 138146 856
rect 138314 575 138422 856
rect 138590 575 138698 856
rect 138866 575 138974 856
rect 139142 575 139342 856
rect 139510 575 139618 856
rect 139786 575 139894 856
rect 140062 575 140262 856
rect 140430 575 140538 856
rect 140706 575 140814 856
rect 140982 575 141182 856
rect 141350 575 141458 856
rect 141626 575 141734 856
rect 141902 575 142102 856
rect 142270 575 142378 856
rect 142546 575 142654 856
rect 142822 575 142930 856
rect 143098 575 143298 856
rect 143466 575 143574 856
rect 143742 575 143850 856
rect 144018 575 144218 856
rect 144386 575 144494 856
rect 144662 575 144770 856
rect 144938 575 145138 856
rect 145306 575 145414 856
rect 145582 575 145690 856
rect 145858 575 146058 856
rect 146226 575 146334 856
rect 146502 575 146610 856
rect 146778 575 146886 856
rect 147054 575 147254 856
rect 147422 575 147530 856
rect 147698 575 147806 856
rect 147974 575 148174 856
rect 148342 575 148450 856
rect 148618 575 148726 856
rect 148894 575 149094 856
rect 149262 575 149370 856
rect 149538 575 149646 856
<< metal3 >>
rect 0 49376 800 49496
rect 149200 49376 150000 49496
rect 0 48152 800 48272
rect 149200 48288 150000 48408
rect 149200 47200 150000 47320
rect 0 46928 800 47048
rect 149200 46112 150000 46232
rect 0 45704 800 45824
rect 149200 45024 150000 45144
rect 0 44616 800 44736
rect 149200 43800 150000 43920
rect 0 43392 800 43512
rect 149200 42712 150000 42832
rect 0 42168 800 42288
rect 149200 41624 150000 41744
rect 0 40944 800 41064
rect 149200 40536 150000 40656
rect 0 39856 800 39976
rect 149200 39448 150000 39568
rect 0 38632 800 38752
rect 149200 38360 150000 38480
rect 0 37408 800 37528
rect 149200 37136 150000 37256
rect 0 36184 800 36304
rect 149200 36048 150000 36168
rect 0 35096 800 35216
rect 149200 34960 150000 35080
rect 0 33872 800 33992
rect 149200 33872 150000 33992
rect 0 32648 800 32768
rect 149200 32784 150000 32904
rect 0 31424 800 31544
rect 149200 31560 150000 31680
rect 0 30336 800 30456
rect 149200 30472 150000 30592
rect 149200 29384 150000 29504
rect 0 29112 800 29232
rect 149200 28296 150000 28416
rect 0 27888 800 28008
rect 149200 27208 150000 27328
rect 0 26664 800 26784
rect 149200 26120 150000 26240
rect 0 25576 800 25696
rect 149200 24896 150000 25016
rect 0 24352 800 24472
rect 149200 23808 150000 23928
rect 0 23128 800 23248
rect 149200 22720 150000 22840
rect 0 21904 800 22024
rect 149200 21632 150000 21752
rect 0 20680 800 20800
rect 149200 20544 150000 20664
rect 0 19592 800 19712
rect 149200 19456 150000 19576
rect 0 18368 800 18488
rect 149200 18232 150000 18352
rect 0 17144 800 17264
rect 149200 17144 150000 17264
rect 0 15920 800 16040
rect 149200 16056 150000 16176
rect 0 14832 800 14952
rect 149200 14968 150000 15088
rect 149200 13880 150000 14000
rect 0 13608 800 13728
rect 149200 12656 150000 12776
rect 0 12384 800 12504
rect 149200 11568 150000 11688
rect 0 11160 800 11280
rect 149200 10480 150000 10600
rect 0 10072 800 10192
rect 149200 9392 150000 9512
rect 0 8848 800 8968
rect 149200 8304 150000 8424
rect 0 7624 800 7744
rect 149200 7216 150000 7336
rect 0 6400 800 6520
rect 149200 5992 150000 6112
rect 0 5312 800 5432
rect 149200 4904 150000 5024
rect 0 4088 800 4208
rect 149200 3816 150000 3936
rect 0 2864 800 2984
rect 149200 2728 150000 2848
rect 0 1640 800 1760
rect 149200 1640 150000 1760
rect 0 552 800 672
rect 149200 552 150000 672
<< obsm3 >>
rect 880 49296 149120 49469
rect 800 48488 149200 49296
rect 800 48352 149120 48488
rect 880 48208 149120 48352
rect 880 48072 149200 48208
rect 800 47400 149200 48072
rect 800 47128 149120 47400
rect 880 47120 149120 47128
rect 880 46848 149200 47120
rect 800 46312 149200 46848
rect 800 46032 149120 46312
rect 800 45904 149200 46032
rect 880 45624 149200 45904
rect 800 45224 149200 45624
rect 800 44944 149120 45224
rect 800 44816 149200 44944
rect 880 44536 149200 44816
rect 800 44000 149200 44536
rect 800 43720 149120 44000
rect 800 43592 149200 43720
rect 880 43312 149200 43592
rect 800 42912 149200 43312
rect 800 42632 149120 42912
rect 800 42368 149200 42632
rect 880 42088 149200 42368
rect 800 41824 149200 42088
rect 800 41544 149120 41824
rect 800 41144 149200 41544
rect 880 40864 149200 41144
rect 800 40736 149200 40864
rect 800 40456 149120 40736
rect 800 40056 149200 40456
rect 880 39776 149200 40056
rect 800 39648 149200 39776
rect 800 39368 149120 39648
rect 800 38832 149200 39368
rect 880 38560 149200 38832
rect 880 38552 149120 38560
rect 800 38280 149120 38552
rect 800 37608 149200 38280
rect 880 37336 149200 37608
rect 880 37328 149120 37336
rect 800 37056 149120 37328
rect 800 36384 149200 37056
rect 880 36248 149200 36384
rect 880 36104 149120 36248
rect 800 35968 149120 36104
rect 800 35296 149200 35968
rect 880 35160 149200 35296
rect 880 35016 149120 35160
rect 800 34880 149120 35016
rect 800 34072 149200 34880
rect 880 33792 149120 34072
rect 800 32984 149200 33792
rect 800 32848 149120 32984
rect 880 32704 149120 32848
rect 880 32568 149200 32704
rect 800 31760 149200 32568
rect 800 31624 149120 31760
rect 880 31480 149120 31624
rect 880 31344 149200 31480
rect 800 30672 149200 31344
rect 800 30536 149120 30672
rect 880 30392 149120 30536
rect 880 30256 149200 30392
rect 800 29584 149200 30256
rect 800 29312 149120 29584
rect 880 29304 149120 29312
rect 880 29032 149200 29304
rect 800 28496 149200 29032
rect 800 28216 149120 28496
rect 800 28088 149200 28216
rect 880 27808 149200 28088
rect 800 27408 149200 27808
rect 800 27128 149120 27408
rect 800 26864 149200 27128
rect 880 26584 149200 26864
rect 800 26320 149200 26584
rect 800 26040 149120 26320
rect 800 25776 149200 26040
rect 880 25496 149200 25776
rect 800 25096 149200 25496
rect 800 24816 149120 25096
rect 800 24552 149200 24816
rect 880 24272 149200 24552
rect 800 24008 149200 24272
rect 800 23728 149120 24008
rect 800 23328 149200 23728
rect 880 23048 149200 23328
rect 800 22920 149200 23048
rect 800 22640 149120 22920
rect 800 22104 149200 22640
rect 880 21832 149200 22104
rect 880 21824 149120 21832
rect 800 21552 149120 21824
rect 800 20880 149200 21552
rect 880 20744 149200 20880
rect 880 20600 149120 20744
rect 800 20464 149120 20600
rect 800 19792 149200 20464
rect 880 19656 149200 19792
rect 880 19512 149120 19656
rect 800 19376 149120 19512
rect 800 18568 149200 19376
rect 880 18432 149200 18568
rect 880 18288 149120 18432
rect 800 18152 149120 18288
rect 800 17344 149200 18152
rect 880 17064 149120 17344
rect 800 16256 149200 17064
rect 800 16120 149120 16256
rect 880 15976 149120 16120
rect 880 15840 149200 15976
rect 800 15168 149200 15840
rect 800 15032 149120 15168
rect 880 14888 149120 15032
rect 880 14752 149200 14888
rect 800 14080 149200 14752
rect 800 13808 149120 14080
rect 880 13800 149120 13808
rect 880 13528 149200 13800
rect 800 12856 149200 13528
rect 800 12584 149120 12856
rect 880 12576 149120 12584
rect 880 12304 149200 12576
rect 800 11768 149200 12304
rect 800 11488 149120 11768
rect 800 11360 149200 11488
rect 880 11080 149200 11360
rect 800 10680 149200 11080
rect 800 10400 149120 10680
rect 800 10272 149200 10400
rect 880 9992 149200 10272
rect 800 9592 149200 9992
rect 800 9312 149120 9592
rect 800 9048 149200 9312
rect 880 8768 149200 9048
rect 800 8504 149200 8768
rect 800 8224 149120 8504
rect 800 7824 149200 8224
rect 880 7544 149200 7824
rect 800 7416 149200 7544
rect 800 7136 149120 7416
rect 800 6600 149200 7136
rect 880 6320 149200 6600
rect 800 6192 149200 6320
rect 800 5912 149120 6192
rect 800 5512 149200 5912
rect 880 5232 149200 5512
rect 800 5104 149200 5232
rect 800 4824 149120 5104
rect 800 4288 149200 4824
rect 880 4016 149200 4288
rect 880 4008 149120 4016
rect 800 3736 149120 4008
rect 800 3064 149200 3736
rect 880 2928 149200 3064
rect 880 2784 149120 2928
rect 800 2648 149120 2784
rect 800 1840 149200 2648
rect 880 1560 149120 1840
rect 800 752 149200 1560
rect 880 579 149120 752
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
rect 65648 2128 65968 47376
rect 81008 2128 81328 47376
rect 96368 2128 96688 47376
rect 111728 2128 112048 47376
rect 127088 2128 127408 47376
rect 142448 2128 142768 47376
<< labels >>
rlabel metal3 s 149200 552 150000 672 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 149200 33872 150000 33992 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 149200 37136 150000 37256 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 149200 40536 150000 40656 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 149200 43800 150000 43920 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 149200 47200 150000 47320 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 147126 49200 147182 50000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 130474 49200 130530 50000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 113822 49200 113878 50000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 97170 49200 97226 50000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 80518 49200 80574 50000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 149200 3816 150000 3936 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 63866 49200 63922 50000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 47122 49200 47178 50000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 30470 49200 30526 50000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 13818 49200 13874 50000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 149200 7216 150000 7336 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 149200 10480 150000 10600 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 149200 13880 150000 14000 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 149200 17144 150000 17264 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 149200 20544 150000 20664 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 149200 23808 150000 23928 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 149200 27208 150000 27328 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 149200 30472 150000 30592 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 149200 2728 150000 2848 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 149200 36048 150000 36168 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 149200 39448 150000 39568 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 149200 42712 150000 42832 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 149200 46112 150000 46232 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 149200 49376 150000 49496 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 135994 49200 136050 50000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 119342 49200 119398 50000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 102690 49200 102746 50000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 86038 49200 86094 50000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 69386 49200 69442 50000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 149200 5992 150000 6112 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 52734 49200 52790 50000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 36082 49200 36138 50000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 19430 49200 19486 50000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 2778 49200 2834 50000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 149200 9392 150000 9512 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 552 800 672 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 149200 12656 150000 12776 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 149200 16056 150000 16176 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 149200 19456 150000 19576 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 149200 22720 150000 22840 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 149200 26120 150000 26240 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 149200 29384 150000 29504 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 149200 32784 150000 32904 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 149200 1640 150000 1760 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 149200 34960 150000 35080 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 149200 38360 150000 38480 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 149200 41624 150000 41744 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 149200 45024 150000 45144 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 149200 48288 150000 48408 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 141606 49200 141662 50000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 124954 49200 125010 50000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 108302 49200 108358 50000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 91558 49200 91614 50000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 74906 49200 74962 50000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 149200 4904 150000 5024 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 58254 49200 58310 50000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 41602 49200 41658 50000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 24950 49200 25006 50000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 8298 49200 8354 50000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 149200 8304 150000 8424 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 149200 11568 150000 11688 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 149200 14968 150000 15088 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 149200 18232 150000 18352 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 149200 21632 150000 21752 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 149200 24896 150000 25016 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 149200 28296 150000 28416 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 149200 31560 150000 31680 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 47376 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 47376 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 47376 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 47376 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 47376 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 47376 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7246388
string GDS_FILE /home/tutel/caravel_tutorial/RNG-SCROLL/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 655732
<< end >>

