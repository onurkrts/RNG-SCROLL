magic
tech sky130A
magscale 1 2
timestamp 1654667515
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 328454 700816 328460 700868
rect 328512 700856 328518 700868
rect 397454 700856 397460 700868
rect 328512 700828 397460 700856
rect 328512 700816 328518 700828
rect 397454 700816 397460 700828
rect 397512 700816 397518 700868
rect 335354 700748 335360 700800
rect 335412 700788 335418 700800
rect 413646 700788 413652 700800
rect 335412 700760 413652 700788
rect 335412 700748 335418 700760
rect 413646 700748 413652 700760
rect 413704 700748 413710 700800
rect 343634 700680 343640 700732
rect 343692 700720 343698 700732
rect 429838 700720 429844 700732
rect 343692 700692 429844 700720
rect 343692 700680 343698 700692
rect 429838 700680 429844 700692
rect 429896 700680 429902 700732
rect 350534 700612 350540 700664
rect 350592 700652 350598 700664
rect 462314 700652 462320 700664
rect 350592 700624 462320 700652
rect 350592 700612 350598 700624
rect 462314 700612 462320 700624
rect 462372 700612 462378 700664
rect 357434 700544 357440 700596
rect 357492 700584 357498 700596
rect 478506 700584 478512 700596
rect 357492 700556 478512 700584
rect 357492 700544 357498 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 365714 700476 365720 700528
rect 365772 700516 365778 700528
rect 494790 700516 494796 700528
rect 365772 700488 494796 700516
rect 365772 700476 365778 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 306374 700408 306380 700460
rect 306432 700448 306438 700460
rect 332502 700448 332508 700460
rect 306432 700420 332508 700448
rect 306432 700408 306438 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 372614 700408 372620 700460
rect 372672 700448 372678 700460
rect 527174 700448 527180 700460
rect 372672 700420 527180 700448
rect 372672 700408 372678 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 313274 700340 313280 700392
rect 313332 700380 313338 700392
rect 348786 700380 348792 700392
rect 313332 700352 348792 700380
rect 313332 700340 313338 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 379514 700340 379520 700392
rect 379572 700380 379578 700392
rect 543458 700380 543464 700392
rect 379572 700352 543464 700380
rect 379572 700340 379578 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 321554 700272 321560 700324
rect 321612 700312 321618 700324
rect 364978 700312 364984 700324
rect 321612 700284 364984 700312
rect 321612 700272 321618 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 387794 700272 387800 700324
rect 387852 700312 387858 700324
rect 559650 700312 559656 700324
rect 387852 700284 559656 700312
rect 387852 700272 387858 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 18598 683176 18604 683188
rect 3476 683148 18604 683176
rect 3476 683136 3482 683148
rect 18598 683136 18604 683148
rect 18656 683136 18662 683188
rect 406378 683136 406384 683188
rect 406436 683176 406442 683188
rect 579614 683176 579620 683188
rect 406436 683148 579620 683176
rect 406436 683136 406442 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 395338 670692 395344 670744
rect 395396 670732 395402 670744
rect 580166 670732 580172 670744
rect 395396 670704 580172 670732
rect 395396 670692 395402 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 400858 643084 400864 643136
rect 400916 643124 400922 643136
rect 580166 643124 580172 643136
rect 400916 643096 580172 643124
rect 400916 643084 400922 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3326 632068 3332 632120
rect 3384 632108 3390 632120
rect 21358 632108 21364 632120
rect 3384 632080 21364 632108
rect 3384 632068 3390 632080
rect 21358 632068 21364 632080
rect 21416 632068 21422 632120
rect 393958 630640 393964 630692
rect 394016 630680 394022 630692
rect 579982 630680 579988 630692
rect 394016 630652 579988 630680
rect 394016 630640 394022 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 13078 618304 13084 618316
rect 3384 618276 13084 618304
rect 3384 618264 3390 618276
rect 13078 618264 13084 618276
rect 13136 618264 13142 618316
rect 2774 605888 2780 605940
rect 2832 605928 2838 605940
rect 4798 605928 4804 605940
rect 2832 605900 4804 605928
rect 2832 605888 2838 605900
rect 4798 605888 4804 605900
rect 4856 605888 4862 605940
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 22738 579680 22744 579692
rect 3384 579652 22744 579680
rect 3384 579640 3390 579652
rect 22738 579640 22744 579652
rect 22796 579640 22802 579692
rect 404998 576852 405004 576904
rect 405056 576892 405062 576904
rect 579982 576892 579988 576904
rect 405056 576864 579988 576892
rect 405056 576852 405062 576864
rect 579982 576852 579988 576864
rect 580040 576852 580046 576904
rect 399478 536800 399484 536852
rect 399536 536840 399542 536852
rect 579614 536840 579620 536852
rect 399536 536812 579620 536840
rect 399536 536800 399542 536812
rect 579614 536800 579620 536812
rect 579672 536800 579678 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 26878 527184 26884 527196
rect 3016 527156 26884 527184
rect 3016 527144 3022 527156
rect 26878 527144 26884 527156
rect 26936 527144 26942 527196
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 14458 514808 14464 514820
rect 3384 514780 14464 514808
rect 3384 514768 3390 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 3326 501304 3332 501356
rect 3384 501344 3390 501356
rect 8938 501344 8944 501356
rect 3384 501316 8944 501344
rect 3384 501304 3390 501316
rect 8938 501304 8944 501316
rect 8996 501304 9002 501356
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 32398 474756 32404 474768
rect 3384 474728 32404 474756
rect 3384 474716 3390 474728
rect 32398 474716 32404 474728
rect 32456 474716 32462 474768
rect 403618 470568 403624 470620
rect 403676 470608 403682 470620
rect 579982 470608 579988 470620
rect 403676 470580 579988 470608
rect 403676 470568 403682 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 549898 456764 549904 456816
rect 549956 456804 549962 456816
rect 580166 456804 580172 456816
rect 549956 456776 580172 456804
rect 549956 456764 549962 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 407758 418140 407764 418192
rect 407816 418180 407822 418192
rect 580166 418180 580172 418192
rect 407816 418152 580172 418180
rect 407816 418140 407822 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 17218 409884 17224 409896
rect 3384 409856 17224 409884
rect 3384 409844 3390 409856
rect 17218 409844 17224 409856
rect 17276 409844 17282 409896
rect 396718 404336 396724 404388
rect 396776 404376 396782 404388
rect 580166 404376 580172 404388
rect 396776 404348 580172 404376
rect 396776 404336 396782 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 10318 397508 10324 397520
rect 3384 397480 10324 397508
rect 3384 397468 3390 397480
rect 10318 397468 10324 397480
rect 10376 397468 10382 397520
rect 169754 393116 169760 393168
rect 169812 393156 169818 393168
rect 254946 393156 254952 393168
rect 169812 393128 254952 393156
rect 169812 393116 169818 393128
rect 254946 393116 254952 393128
rect 255004 393116 255010 393168
rect 153194 393048 153200 393100
rect 153252 393088 153258 393100
rect 247494 393088 247500 393100
rect 153252 393060 247500 393088
rect 153252 393048 153258 393060
rect 247494 393048 247500 393060
rect 247552 393048 247558 393100
rect 136634 392980 136640 393032
rect 136692 393020 136698 393032
rect 240134 393020 240140 393032
rect 136692 392992 240140 393020
rect 136692 392980 136698 392992
rect 240134 392980 240140 392992
rect 240192 392980 240198 393032
rect 104894 392912 104900 392964
rect 104952 392952 104958 392964
rect 232682 392952 232688 392964
rect 104952 392924 232688 392952
rect 104952 392912 104958 392924
rect 232682 392912 232688 392924
rect 232740 392912 232746 392964
rect 88334 392844 88340 392896
rect 88392 392884 88398 392896
rect 225322 392884 225328 392896
rect 88392 392856 225328 392884
rect 88392 392844 88398 392856
rect 225322 392844 225328 392856
rect 225380 392844 225386 392896
rect 71774 392776 71780 392828
rect 71832 392816 71838 392828
rect 217870 392816 217876 392828
rect 71832 392788 217876 392816
rect 71832 392776 71838 392788
rect 217870 392776 217876 392788
rect 217928 392776 217934 392828
rect 40034 392708 40040 392760
rect 40092 392748 40098 392760
rect 210510 392748 210516 392760
rect 40092 392720 210516 392748
rect 40092 392708 40098 392720
rect 210510 392708 210516 392720
rect 210568 392708 210574 392760
rect 234614 392708 234620 392760
rect 234672 392748 234678 392760
rect 277118 392748 277124 392760
rect 234672 392720 277124 392748
rect 234672 392708 234678 392720
rect 277118 392708 277124 392720
rect 277176 392708 277182 392760
rect 23474 392640 23480 392692
rect 23532 392680 23538 392692
rect 203058 392680 203064 392692
rect 23532 392652 203064 392680
rect 23532 392640 23538 392652
rect 203058 392640 203064 392652
rect 203116 392640 203122 392692
rect 218054 392640 218060 392692
rect 218112 392680 218118 392692
rect 269758 392680 269764 392692
rect 218112 392652 269764 392680
rect 218112 392640 218118 392652
rect 269758 392640 269764 392652
rect 269816 392640 269822 392692
rect 282914 392640 282920 392692
rect 282972 392680 282978 392692
rect 291930 392680 291936 392692
rect 282972 392652 291936 392680
rect 282972 392640 282978 392652
rect 291930 392640 291936 392652
rect 291988 392640 291994 392692
rect 6914 392572 6920 392624
rect 6972 392612 6978 392624
rect 195698 392612 195704 392624
rect 6972 392584 195704 392612
rect 6972 392572 6978 392584
rect 195698 392572 195704 392584
rect 195756 392572 195762 392624
rect 201494 392572 201500 392624
rect 201552 392612 201558 392624
rect 262306 392612 262312 392624
rect 201552 392584 262312 392612
rect 201552 392572 201558 392584
rect 262306 392572 262312 392584
rect 262364 392572 262370 392624
rect 266354 392572 266360 392624
rect 266412 392612 266418 392624
rect 284570 392612 284576 392624
rect 266412 392584 284576 392612
rect 266412 392572 266418 392584
rect 284570 392572 284576 392584
rect 284628 392572 284634 392624
rect 18598 387744 18604 387796
rect 18656 387784 18662 387796
rect 189074 387784 189080 387796
rect 18656 387756 189080 387784
rect 18656 387744 18662 387756
rect 189074 387744 189080 387756
rect 189132 387744 189138 387796
rect 394510 387744 394516 387796
rect 394568 387784 394574 387796
rect 580258 387784 580264 387796
rect 394568 387756 580264 387784
rect 394568 387744 394574 387756
rect 580258 387744 580264 387756
rect 580316 387744 580322 387796
rect 3418 380808 3424 380860
rect 3476 380848 3482 380860
rect 189074 380848 189080 380860
rect 3476 380820 189080 380848
rect 3476 380808 3482 380820
rect 189074 380808 189080 380820
rect 189132 380808 189138 380860
rect 394602 380808 394608 380860
rect 394660 380848 394666 380860
rect 406378 380848 406384 380860
rect 394660 380820 406384 380848
rect 394660 380808 394666 380820
rect 406378 380808 406384 380820
rect 406436 380808 406442 380860
rect 394142 375300 394148 375352
rect 394200 375340 394206 375352
rect 395338 375340 395344 375352
rect 394200 375312 395344 375340
rect 394200 375300 394206 375312
rect 395338 375300 395344 375312
rect 395396 375300 395402 375352
rect 3510 373940 3516 373992
rect 3568 373980 3574 373992
rect 189074 373980 189080 373992
rect 3568 373952 189080 373980
rect 3568 373940 3574 373952
rect 189074 373940 189080 373952
rect 189132 373940 189138 373992
rect 393866 368092 393872 368144
rect 393924 368132 393930 368144
rect 400858 368132 400864 368144
rect 393924 368104 400864 368132
rect 393924 368092 393930 368104
rect 400858 368092 400864 368104
rect 400916 368092 400922 368144
rect 21358 367004 21364 367056
rect 21416 367044 21422 367056
rect 189074 367044 189080 367056
rect 21416 367016 189080 367044
rect 21416 367004 21422 367016
rect 189074 367004 189080 367016
rect 189132 367004 189138 367056
rect 394050 364352 394056 364404
rect 394108 364392 394114 364404
rect 580166 364392 580172 364404
rect 394108 364364 580172 364392
rect 394108 364352 394114 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 13078 360136 13084 360188
rect 13136 360176 13142 360188
rect 189074 360176 189080 360188
rect 13136 360148 189080 360176
rect 13136 360136 13142 360148
rect 189074 360136 189080 360148
rect 189132 360136 189138 360188
rect 394602 355988 394608 356040
rect 394660 356028 394666 356040
rect 580350 356028 580356 356040
rect 394660 356000 580356 356028
rect 394660 355988 394666 356000
rect 580350 355988 580356 356000
rect 580408 355988 580414 356040
rect 4798 353200 4804 353252
rect 4856 353240 4862 353252
rect 189074 353240 189080 353252
rect 4856 353212 189080 353240
rect 4856 353200 4862 353212
rect 189074 353200 189080 353212
rect 189132 353200 189138 353252
rect 394602 350480 394608 350532
rect 394660 350520 394666 350532
rect 580442 350520 580448 350532
rect 394660 350492 580448 350520
rect 394660 350480 394666 350492
rect 580442 350480 580448 350492
rect 580500 350480 580506 350532
rect 22738 347692 22744 347744
rect 22796 347732 22802 347744
rect 189074 347732 189080 347744
rect 22796 347704 189080 347732
rect 22796 347692 22802 347704
rect 189074 347692 189080 347704
rect 189132 347692 189138 347744
rect 394234 343544 394240 343596
rect 394292 343584 394298 343596
rect 404998 343584 405004 343596
rect 394292 343556 405004 343584
rect 394292 343544 394298 343556
rect 404998 343544 405004 343556
rect 405056 343544 405062 343596
rect 3602 340824 3608 340876
rect 3660 340864 3666 340876
rect 189074 340864 189080 340876
rect 3660 340836 189080 340864
rect 3660 340824 3666 340836
rect 189074 340824 189080 340836
rect 189132 340824 189138 340876
rect 394602 338036 394608 338088
rect 394660 338076 394666 338088
rect 580534 338076 580540 338088
rect 394660 338048 580540 338076
rect 394660 338036 394666 338048
rect 580534 338036 580540 338048
rect 580592 338036 580598 338088
rect 3694 333888 3700 333940
rect 3752 333928 3758 333940
rect 189074 333928 189080 333940
rect 3752 333900 189080 333928
rect 3752 333888 3758 333900
rect 189074 333888 189080 333900
rect 189132 333888 189138 333940
rect 393958 331168 393964 331220
rect 394016 331208 394022 331220
rect 399478 331208 399484 331220
rect 394016 331180 399484 331208
rect 394016 331168 394022 331180
rect 399478 331168 399484 331180
rect 399536 331168 399542 331220
rect 26878 327020 26884 327072
rect 26936 327060 26942 327072
rect 189074 327060 189080 327072
rect 26936 327032 189080 327060
rect 26936 327020 26942 327032
rect 189074 327020 189080 327032
rect 189132 327020 189138 327072
rect 394602 325592 394608 325644
rect 394660 325632 394666 325644
rect 580626 325632 580632 325644
rect 394660 325604 580632 325632
rect 394660 325592 394666 325604
rect 580626 325592 580632 325604
rect 580684 325592 580690 325644
rect 14458 320084 14464 320136
rect 14516 320124 14522 320136
rect 189074 320124 189080 320136
rect 14516 320096 189080 320124
rect 14516 320084 14522 320096
rect 189074 320084 189080 320096
rect 189132 320084 189138 320136
rect 394602 318724 394608 318776
rect 394660 318764 394666 318776
rect 580718 318764 580724 318776
rect 394660 318736 580724 318764
rect 394660 318724 394666 318736
rect 580718 318724 580724 318736
rect 580776 318724 580782 318776
rect 8938 314576 8944 314628
rect 8996 314616 9002 314628
rect 189074 314616 189080 314628
rect 8996 314588 189080 314616
rect 8996 314576 9002 314588
rect 189074 314576 189080 314588
rect 189132 314576 189138 314628
rect 394602 313216 394608 313268
rect 394660 313256 394666 313268
rect 580810 313256 580816 313268
rect 394660 313228 580816 313256
rect 394660 313216 394666 313228
rect 580810 313216 580816 313228
rect 580868 313216 580874 313268
rect 393958 311856 393964 311908
rect 394016 311896 394022 311908
rect 580166 311896 580172 311908
rect 394016 311868 580172 311896
rect 394016 311856 394022 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 32398 307708 32404 307760
rect 32456 307748 32462 307760
rect 189074 307748 189080 307760
rect 32456 307720 189080 307748
rect 32456 307708 32462 307720
rect 189074 307708 189080 307720
rect 189132 307708 189138 307760
rect 394234 306280 394240 306332
rect 394292 306320 394298 306332
rect 403618 306320 403624 306332
rect 394292 306292 403624 306320
rect 394292 306280 394298 306292
rect 403618 306280 403624 306292
rect 403676 306280 403682 306332
rect 3786 300772 3792 300824
rect 3844 300812 3850 300824
rect 189074 300812 189080 300824
rect 3844 300784 189080 300812
rect 3844 300772 3850 300784
rect 189074 300772 189080 300784
rect 189132 300772 189138 300824
rect 394602 300772 394608 300824
rect 394660 300812 394666 300824
rect 549898 300812 549904 300824
rect 394660 300784 549904 300812
rect 394660 300772 394666 300784
rect 549898 300772 549904 300784
rect 549956 300772 549962 300824
rect 3878 293904 3884 293956
rect 3936 293944 3942 293956
rect 189074 293944 189080 293956
rect 3936 293916 189080 293944
rect 3936 293904 3942 293916
rect 189074 293904 189080 293916
rect 189132 293904 189138 293956
rect 394602 293904 394608 293956
rect 394660 293944 394666 293956
rect 580902 293944 580908 293956
rect 394660 293916 580908 293944
rect 394660 293904 394666 293916
rect 580902 293904 580908 293916
rect 580960 293904 580966 293956
rect 394602 288328 394608 288380
rect 394660 288368 394666 288380
rect 407758 288368 407764 288380
rect 394660 288340 407764 288368
rect 394660 288328 394666 288340
rect 407758 288328 407764 288340
rect 407816 288328 407822 288380
rect 3970 286968 3976 287020
rect 4028 287008 4034 287020
rect 189074 287008 189080 287020
rect 4028 286980 189080 287008
rect 4028 286968 4034 286980
rect 189074 286968 189080 286980
rect 189132 286968 189138 287020
rect 393682 281256 393688 281308
rect 393740 281296 393746 281308
rect 396718 281296 396724 281308
rect 393740 281268 396724 281296
rect 393740 281256 393746 281268
rect 396718 281256 396724 281268
rect 396776 281256 396782 281308
rect 17218 280100 17224 280152
rect 17276 280140 17282 280152
rect 189074 280140 189080 280152
rect 17276 280112 189080 280140
rect 17276 280100 17282 280112
rect 189074 280100 189080 280112
rect 189132 280100 189138 280152
rect 394602 275952 394608 276004
rect 394660 275992 394666 276004
rect 580258 275992 580264 276004
rect 394660 275964 580264 275992
rect 394660 275952 394666 275964
rect 580258 275952 580264 275964
rect 580316 275952 580322 276004
rect 10318 274592 10324 274644
rect 10376 274632 10382 274644
rect 189074 274632 189080 274644
rect 10376 274604 189080 274632
rect 10376 274592 10382 274604
rect 189074 274592 189080 274604
rect 189132 274592 189138 274644
rect 3418 267656 3424 267708
rect 3476 267696 3482 267708
rect 189074 267696 189080 267708
rect 3476 267668 189080 267696
rect 3476 267656 3482 267668
rect 189074 267656 189080 267668
rect 189132 267656 189138 267708
rect 394602 263508 394608 263560
rect 394660 263548 394666 263560
rect 580350 263548 580356 263560
rect 394660 263520 580356 263548
rect 394660 263508 394666 263520
rect 580350 263508 580356 263520
rect 580408 263508 580414 263560
rect 3510 260788 3516 260840
rect 3568 260828 3574 260840
rect 189074 260828 189080 260840
rect 3568 260800 189080 260828
rect 3568 260788 3574 260800
rect 189074 260788 189080 260800
rect 189132 260788 189138 260840
rect 394050 258068 394056 258120
rect 394108 258108 394114 258120
rect 580166 258108 580172 258120
rect 394108 258080 580172 258108
rect 394108 258068 394114 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 394602 256640 394608 256692
rect 394660 256680 394666 256692
rect 580442 256680 580448 256692
rect 394660 256652 580448 256680
rect 394660 256640 394666 256652
rect 580442 256640 580448 256652
rect 580500 256640 580506 256692
rect 4062 253852 4068 253904
rect 4120 253892 4126 253904
rect 189074 253892 189080 253904
rect 4120 253864 189080 253892
rect 4120 253852 4126 253864
rect 189074 253852 189080 253864
rect 189132 253852 189138 253904
rect 3602 246984 3608 247036
rect 3660 247024 3666 247036
rect 189074 247024 189080 247036
rect 3660 246996 189080 247024
rect 3660 246984 3666 246996
rect 189074 246984 189080 246996
rect 189132 246984 189138 247036
rect 394602 244196 394608 244248
rect 394660 244236 394666 244248
rect 580534 244236 580540 244248
rect 394660 244208 580540 244236
rect 394660 244196 394666 244208
rect 580534 244196 580540 244208
rect 580592 244196 580598 244248
rect 3694 240048 3700 240100
rect 3752 240088 3758 240100
rect 189074 240088 189080 240100
rect 3752 240060 189080 240088
rect 3752 240048 3758 240060
rect 189074 240048 189080 240060
rect 189132 240048 189138 240100
rect 394602 238688 394608 238740
rect 394660 238728 394666 238740
rect 580258 238728 580264 238740
rect 394660 238700 580264 238728
rect 394660 238688 394666 238700
rect 580258 238688 580264 238700
rect 580316 238688 580322 238740
rect 3786 234540 3792 234592
rect 3844 234580 3850 234592
rect 189074 234580 189080 234592
rect 3844 234552 189080 234580
rect 3844 234540 3850 234552
rect 189074 234540 189080 234552
rect 189132 234540 189138 234592
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 579798 231860 579804 231872
rect 394016 231832 579804 231860
rect 394016 231820 394022 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 3878 227672 3884 227724
rect 3936 227712 3942 227724
rect 189074 227712 189080 227724
rect 3936 227684 189080 227712
rect 3936 227672 3942 227684
rect 189074 227672 189080 227684
rect 189132 227672 189138 227724
rect 394602 226244 394608 226296
rect 394660 226284 394666 226296
rect 580350 226284 580356 226296
rect 394660 226256 580356 226284
rect 394660 226244 394666 226256
rect 580350 226244 580356 226256
rect 580408 226244 580414 226296
rect 3418 220736 3424 220788
rect 3476 220776 3482 220788
rect 189074 220776 189080 220788
rect 3476 220748 189080 220776
rect 3476 220736 3482 220748
rect 189074 220736 189080 220748
rect 189132 220736 189138 220788
rect 393958 218016 393964 218068
rect 394016 218056 394022 218068
rect 580166 218056 580172 218068
rect 394016 218028 580172 218056
rect 394016 218016 394022 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3510 213868 3516 213920
rect 3568 213908 3574 213920
rect 189074 213908 189080 213920
rect 3568 213880 189080 213908
rect 3568 213868 3574 213880
rect 189074 213868 189080 213880
rect 189132 213868 189138 213920
rect 3418 206932 3424 206984
rect 3476 206972 3482 206984
rect 189074 206972 189080 206984
rect 3476 206944 189080 206972
rect 3476 206932 3482 206944
rect 189074 206932 189080 206944
rect 189132 206932 189138 206984
rect 394602 206252 394608 206304
rect 394660 206292 394666 206304
rect 580166 206292 580172 206304
rect 394660 206264 580172 206292
rect 394660 206252 394666 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 3142 200064 3148 200116
rect 3200 200104 3206 200116
rect 189074 200104 189080 200116
rect 3200 200076 189080 200104
rect 3200 200064 3206 200076
rect 189074 200064 189080 200076
rect 189132 200064 189138 200116
rect 3418 193196 3424 193248
rect 3476 193236 3482 193248
rect 189074 193236 189080 193248
rect 3476 193208 189080 193236
rect 3476 193196 3482 193208
rect 189074 193196 189080 193208
rect 189132 193196 189138 193248
rect 394050 193128 394056 193180
rect 394108 193168 394114 193180
rect 580166 193168 580172 193180
rect 394108 193140 580172 193168
rect 394108 193128 394114 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3418 179392 3424 179444
rect 3476 179432 3482 179444
rect 189074 179432 189080 179444
rect 3476 179404 189080 179432
rect 3476 179392 3482 179404
rect 189074 179392 189080 179404
rect 189132 179392 189138 179444
rect 393958 179324 393964 179376
rect 394016 179364 394022 179376
rect 580166 179364 580172 179376
rect 394016 179336 580172 179364
rect 394016 179324 394022 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 394234 166948 394240 167000
rect 394292 166988 394298 167000
rect 580166 166988 580172 167000
rect 394292 166960 580172 166988
rect 394292 166948 394298 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 189810 164200 189816 164212
rect 3292 164172 189816 164200
rect 3292 164160 3298 164172
rect 189810 164160 189816 164172
rect 189868 164160 189874 164212
rect 3602 158720 3608 158772
rect 3660 158760 3666 158772
rect 189074 158760 189080 158772
rect 3660 158732 189080 158760
rect 3660 158720 3666 158732
rect 189074 158720 189080 158732
rect 189132 158720 189138 158772
rect 394142 153144 394148 153196
rect 394200 153184 394206 153196
rect 580166 153184 580172 153196
rect 394200 153156 580172 153184
rect 394200 153144 394206 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3510 139408 3516 139460
rect 3568 139448 3574 139460
rect 189074 139448 189080 139460
rect 3568 139420 189080 139448
rect 3568 139408 3574 139420
rect 189074 139408 189080 139420
rect 189132 139408 189138 139460
rect 394050 139340 394056 139392
rect 394108 139380 394114 139392
rect 580166 139380 580172 139392
rect 394108 139352 580172 139380
rect 394108 139340 394114 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3418 137912 3424 137964
rect 3476 137952 3482 137964
rect 189718 137952 189724 137964
rect 3476 137924 189724 137952
rect 3476 137912 3482 137924
rect 189718 137912 189724 137924
rect 189776 137912 189782 137964
rect 393774 131112 393780 131164
rect 393832 131152 393838 131164
rect 395338 131152 395344 131164
rect 393832 131124 395344 131152
rect 393832 131112 393838 131124
rect 395338 131112 395344 131124
rect 395396 131112 395402 131164
rect 393958 126896 393964 126948
rect 394016 126936 394022 126948
rect 580166 126936 580172 126948
rect 394016 126908 580172 126936
rect 394016 126896 394022 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3418 118668 3424 118720
rect 3476 118708 3482 118720
rect 189074 118708 189080 118720
rect 3476 118680 189080 118708
rect 3476 118668 3482 118680
rect 189074 118668 189080 118680
rect 189132 118668 189138 118720
rect 395338 115200 395344 115252
rect 395396 115240 395402 115252
rect 580258 115240 580264 115252
rect 395396 115212 580264 115240
rect 395396 115200 395402 115212
rect 580258 115200 580264 115212
rect 580316 115200 580322 115252
rect 394510 113092 394516 113144
rect 394568 113132 394574 113144
rect 580166 113132 580172 113144
rect 394568 113104 580172 113132
rect 394568 113092 394574 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 394602 111800 394608 111852
rect 394660 111840 394666 111852
rect 395338 111840 395344 111852
rect 394660 111812 395344 111840
rect 394660 111800 394666 111812
rect 395338 111800 395344 111812
rect 395396 111800 395402 111852
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 190178 111772 190184 111784
rect 3384 111744 190184 111772
rect 3384 111732 3390 111744
rect 190178 111732 190184 111744
rect 190236 111732 190242 111784
rect 224954 110168 224960 110220
rect 225012 110208 225018 110220
rect 225138 110208 225144 110220
rect 225012 110180 225144 110208
rect 225012 110168 225018 110180
rect 225138 110168 225144 110180
rect 225196 110168 225202 110220
rect 238754 110168 238760 110220
rect 238812 110208 238818 110220
rect 238938 110208 238944 110220
rect 238812 110180 238944 110208
rect 238812 110168 238818 110180
rect 238938 110168 238944 110180
rect 238996 110168 239002 110220
rect 345014 110168 345020 110220
rect 345072 110208 345078 110220
rect 345198 110208 345204 110220
rect 345072 110180 345204 110208
rect 345072 110168 345078 110180
rect 345198 110168 345204 110180
rect 345256 110168 345262 110220
rect 285674 108808 285680 108860
rect 285732 108848 285738 108860
rect 286318 108848 286324 108860
rect 285732 108820 286324 108848
rect 285732 108808 285738 108820
rect 286318 108808 286324 108820
rect 286376 108808 286382 108860
rect 314654 108808 314660 108860
rect 314712 108848 314718 108860
rect 314838 108848 314844 108860
rect 314712 108820 314844 108848
rect 314712 108808 314718 108820
rect 314838 108808 314844 108820
rect 314896 108808 314902 108860
rect 390554 108672 390560 108724
rect 390612 108712 390618 108724
rect 400858 108712 400864 108724
rect 390612 108684 400864 108712
rect 390612 108672 390618 108684
rect 400858 108672 400864 108684
rect 400916 108672 400922 108724
rect 188338 108604 188344 108656
rect 188396 108644 188402 108656
rect 209590 108644 209596 108656
rect 188396 108616 209596 108644
rect 188396 108604 188402 108616
rect 209590 108604 209596 108616
rect 209648 108604 209654 108656
rect 339402 108604 339408 108656
rect 339460 108644 339466 108656
rect 339460 108616 345014 108644
rect 339460 108604 339466 108616
rect 124214 108536 124220 108588
rect 124272 108576 124278 108588
rect 234798 108576 234804 108588
rect 124272 108548 234804 108576
rect 124272 108536 124278 108548
rect 234798 108536 234804 108548
rect 234856 108536 234862 108588
rect 253198 108536 253204 108588
rect 253256 108576 253262 108588
rect 262306 108576 262312 108588
rect 253256 108548 262312 108576
rect 253256 108536 253262 108548
rect 262306 108536 262312 108548
rect 262364 108536 262370 108588
rect 285950 108536 285956 108588
rect 286008 108576 286014 108588
rect 290366 108576 290372 108588
rect 286008 108548 290372 108576
rect 286008 108536 286014 108548
rect 290366 108536 290372 108548
rect 290424 108536 290430 108588
rect 313090 108536 313096 108588
rect 313148 108576 313154 108588
rect 313148 108548 340184 108576
rect 313148 108536 313154 108548
rect 117314 108468 117320 108520
rect 117372 108508 117378 108520
rect 232314 108508 232320 108520
rect 117372 108480 232320 108508
rect 117372 108468 117378 108480
rect 232314 108468 232320 108480
rect 232372 108468 232378 108520
rect 235350 108468 235356 108520
rect 235408 108508 235414 108520
rect 249794 108508 249800 108520
rect 235408 108480 249800 108508
rect 235408 108468 235414 108480
rect 249794 108468 249800 108480
rect 249852 108468 249858 108520
rect 250438 108468 250444 108520
rect 250496 108508 250502 108520
rect 264330 108508 264336 108520
rect 250496 108480 264336 108508
rect 250496 108468 250502 108480
rect 264330 108468 264336 108480
rect 264388 108468 264394 108520
rect 278774 108468 278780 108520
rect 278832 108508 278838 108520
rect 287882 108508 287888 108520
rect 278832 108480 287888 108508
rect 278832 108468 278838 108480
rect 287882 108468 287888 108480
rect 287940 108468 287946 108520
rect 110414 108400 110420 108452
rect 110472 108440 110478 108452
rect 229922 108440 229928 108452
rect 110472 108412 229928 108440
rect 110472 108400 110478 108412
rect 229922 108400 229928 108412
rect 229980 108400 229986 108452
rect 247678 108400 247684 108452
rect 247736 108440 247742 108452
rect 263134 108440 263140 108452
rect 247736 108412 263140 108440
rect 247736 108400 247742 108412
rect 263134 108400 263140 108412
rect 263192 108400 263198 108452
rect 265618 108400 265624 108452
rect 265676 108440 265682 108452
rect 273806 108440 273812 108452
rect 265676 108412 273812 108440
rect 265676 108400 265682 108412
rect 273806 108400 273812 108412
rect 273864 108400 273870 108452
rect 273898 108400 273904 108452
rect 273956 108440 273962 108452
rect 280154 108440 280160 108452
rect 273956 108412 280160 108440
rect 273956 108400 273962 108412
rect 280154 108400 280160 108412
rect 280212 108400 280218 108452
rect 281534 108400 281540 108452
rect 281592 108440 281598 108452
rect 288710 108440 288716 108452
rect 281592 108412 288716 108440
rect 281592 108400 281598 108412
rect 288710 108400 288716 108412
rect 288768 108400 288774 108452
rect 302878 108400 302884 108452
rect 302936 108440 302942 108452
rect 315298 108440 315304 108452
rect 302936 108412 315304 108440
rect 302936 108400 302942 108412
rect 315298 108400 315304 108412
rect 315356 108400 315362 108452
rect 333330 108400 333336 108452
rect 333388 108440 333394 108452
rect 338666 108440 338672 108452
rect 333388 108412 338672 108440
rect 333388 108400 333394 108412
rect 338666 108400 338672 108412
rect 338724 108400 338730 108452
rect 17218 108332 17224 108384
rect 17276 108372 17282 108384
rect 197446 108372 197452 108384
rect 17276 108344 197452 108372
rect 17276 108332 17282 108344
rect 197446 108332 197452 108344
rect 197504 108332 197510 108384
rect 235258 108332 235264 108384
rect 235316 108372 235322 108384
rect 266814 108372 266820 108384
rect 235316 108344 266820 108372
rect 235316 108332 235322 108344
rect 266814 108332 266820 108344
rect 266872 108332 266878 108384
rect 277762 108332 277768 108384
rect 277820 108372 277826 108384
rect 287514 108372 287520 108384
rect 277820 108344 287520 108372
rect 277820 108332 277826 108344
rect 287514 108332 287520 108344
rect 287572 108332 287578 108384
rect 300026 108332 300032 108384
rect 300084 108372 300090 108384
rect 309778 108372 309784 108384
rect 300084 108344 309784 108372
rect 300084 108332 300090 108344
rect 309778 108332 309784 108344
rect 309836 108332 309842 108384
rect 310606 108332 310612 108384
rect 310664 108372 310670 108384
rect 333238 108372 333244 108384
rect 310664 108344 333244 108372
rect 310664 108332 310670 108344
rect 333238 108332 333244 108344
rect 333296 108332 333302 108384
rect 10318 108264 10324 108316
rect 10376 108304 10382 108316
rect 194226 108304 194232 108316
rect 10376 108276 194232 108304
rect 10376 108264 10382 108276
rect 194226 108264 194232 108276
rect 194284 108264 194290 108316
rect 218698 108264 218704 108316
rect 218756 108304 218762 108316
rect 222194 108304 222200 108316
rect 218756 108276 222200 108304
rect 218756 108264 218762 108276
rect 222194 108264 222200 108276
rect 222252 108264 222258 108316
rect 223574 108264 223580 108316
rect 223632 108304 223638 108316
rect 268838 108304 268844 108316
rect 223632 108276 268844 108304
rect 223632 108264 223638 108276
rect 268838 108264 268844 108276
rect 268896 108264 268902 108316
rect 274634 108264 274640 108316
rect 274692 108304 274698 108316
rect 285674 108304 285680 108316
rect 274692 108276 285680 108304
rect 274692 108264 274698 108276
rect 285674 108264 285680 108276
rect 285732 108264 285738 108316
rect 304902 108264 304908 108316
rect 304960 108304 304966 108316
rect 328454 108304 328460 108316
rect 304960 108276 328460 108304
rect 304960 108264 304966 108276
rect 328454 108264 328460 108276
rect 328512 108264 328518 108316
rect 340156 108304 340184 108548
rect 344986 108508 345014 108616
rect 381170 108604 381176 108656
rect 381228 108644 381234 108656
rect 396718 108644 396724 108656
rect 381228 108616 396724 108644
rect 381228 108604 381234 108616
rect 396718 108604 396724 108616
rect 396776 108604 396782 108656
rect 370222 108536 370228 108588
rect 370280 108576 370286 108588
rect 392578 108576 392584 108588
rect 370280 108548 392584 108576
rect 370280 108536 370286 108548
rect 392578 108536 392584 108548
rect 392636 108536 392642 108588
rect 429194 108508 429200 108520
rect 344986 108480 429200 108508
rect 429194 108468 429200 108480
rect 429252 108468 429258 108520
rect 341886 108400 341892 108452
rect 341944 108440 341950 108452
rect 436094 108440 436100 108452
rect 341944 108412 436100 108440
rect 341944 108400 341950 108412
rect 436094 108400 436100 108412
rect 436152 108400 436158 108452
rect 344278 108332 344284 108384
rect 344336 108372 344342 108384
rect 442994 108372 443000 108384
rect 344336 108344 443000 108372
rect 344336 108332 344342 108344
rect 442994 108332 443000 108344
rect 443052 108332 443058 108384
rect 340156 108276 345014 108304
rect 247218 108128 247224 108180
rect 247276 108168 247282 108180
rect 248506 108168 248512 108180
rect 247276 108140 248512 108168
rect 247276 108128 247282 108140
rect 248506 108128 248512 108140
rect 248564 108128 248570 108180
rect 257430 108128 257436 108180
rect 257488 108168 257494 108180
rect 258258 108168 258264 108180
rect 257488 108140 258264 108168
rect 257488 108128 257494 108140
rect 258258 108128 258264 108140
rect 258316 108128 258322 108180
rect 296714 108128 296720 108180
rect 296772 108168 296778 108180
rect 297358 108168 297364 108180
rect 296772 108140 297364 108168
rect 296772 108128 296778 108140
rect 297358 108128 297364 108140
rect 297416 108128 297422 108180
rect 257338 108060 257344 108112
rect 257396 108100 257402 108112
rect 259086 108100 259092 108112
rect 257396 108072 259092 108100
rect 257396 108060 257402 108072
rect 259086 108060 259092 108072
rect 259144 108060 259150 108112
rect 330110 108060 330116 108112
rect 330168 108100 330174 108112
rect 337378 108100 337384 108112
rect 330168 108072 337384 108100
rect 330168 108060 330174 108072
rect 337378 108060 337384 108072
rect 337436 108060 337442 108112
rect 344986 108100 345014 108276
rect 346762 108264 346768 108316
rect 346820 108304 346826 108316
rect 449894 108304 449900 108316
rect 346820 108276 449900 108304
rect 346820 108264 346826 108276
rect 449894 108264 449900 108276
rect 449952 108264 449958 108316
rect 347038 108100 347044 108112
rect 344986 108072 347044 108100
rect 347038 108060 347044 108072
rect 347096 108060 347102 108112
rect 252002 107992 252008 108044
rect 252060 108032 252066 108044
rect 259546 108032 259552 108044
rect 252060 108004 259552 108032
rect 252060 107992 252066 108004
rect 259546 107992 259552 108004
rect 259604 107992 259610 108044
rect 295242 107992 295248 108044
rect 295300 108032 295306 108044
rect 297358 108032 297364 108044
rect 295300 108004 297364 108032
rect 295300 107992 295306 108004
rect 297358 107992 297364 108004
rect 297416 107992 297422 108044
rect 319990 107924 319996 107976
rect 320048 107964 320054 107976
rect 327626 107964 327632 107976
rect 320048 107936 327632 107964
rect 320048 107924 320054 107936
rect 327626 107924 327632 107936
rect 327684 107924 327690 107976
rect 238110 107788 238116 107840
rect 238168 107828 238174 107840
rect 241238 107828 241244 107840
rect 238168 107800 241244 107828
rect 238168 107788 238174 107800
rect 241238 107788 241244 107800
rect 241296 107788 241302 107840
rect 287422 107788 287428 107840
rect 287480 107828 287486 107840
rect 290734 107828 290740 107840
rect 287480 107800 290740 107828
rect 287480 107788 287486 107800
rect 290734 107788 290740 107800
rect 290792 107788 290798 107840
rect 193858 107720 193864 107772
rect 193916 107760 193922 107772
rect 194962 107760 194968 107772
rect 193916 107732 194968 107760
rect 193916 107720 193922 107732
rect 194962 107720 194968 107732
rect 195020 107720 195026 107772
rect 203518 107720 203524 107772
rect 203576 107760 203582 107772
rect 205174 107760 205180 107772
rect 203576 107732 205180 107760
rect 203576 107720 203582 107732
rect 205174 107720 205180 107732
rect 205232 107720 205238 107772
rect 220078 107720 220084 107772
rect 220136 107760 220142 107772
rect 226610 107760 226616 107772
rect 220136 107732 226616 107760
rect 220136 107720 220142 107732
rect 226610 107720 226616 107732
rect 226668 107720 226674 107772
rect 238018 107720 238024 107772
rect 238076 107760 238082 107772
rect 240410 107760 240416 107772
rect 238076 107732 240416 107760
rect 238076 107720 238082 107732
rect 240410 107720 240416 107732
rect 240468 107720 240474 107772
rect 288434 107720 288440 107772
rect 288492 107760 288498 107772
rect 291102 107760 291108 107772
rect 288492 107732 291108 107760
rect 288492 107720 288498 107732
rect 291102 107720 291108 107732
rect 291160 107720 291166 107772
rect 298462 107720 298468 107772
rect 298520 107760 298526 107772
rect 302878 107760 302884 107772
rect 298520 107732 302884 107760
rect 298520 107720 298526 107732
rect 302878 107720 302884 107732
rect 302936 107720 302942 107772
rect 308582 107720 308588 107772
rect 308640 107760 308646 107772
rect 311250 107760 311256 107772
rect 308640 107732 311256 107760
rect 308640 107720 308646 107732
rect 311250 107720 311256 107732
rect 311308 107720 311314 107772
rect 365806 107720 365812 107772
rect 365864 107760 365870 107772
rect 369118 107760 369124 107772
rect 365864 107732 369124 107760
rect 365864 107720 365870 107732
rect 369118 107720 369124 107732
rect 369176 107720 369182 107772
rect 383654 107720 383660 107772
rect 383712 107760 383718 107772
rect 385862 107760 385868 107772
rect 383712 107732 385868 107760
rect 383712 107720 383718 107732
rect 385862 107720 385868 107732
rect 385920 107720 385926 107772
rect 193950 107652 193956 107704
rect 194008 107692 194014 107704
rect 194594 107692 194600 107704
rect 194008 107664 194600 107692
rect 194008 107652 194014 107664
rect 194594 107652 194600 107664
rect 194652 107652 194658 107704
rect 203702 107652 203708 107704
rect 203760 107692 203766 107704
rect 204714 107692 204720 107704
rect 203760 107664 204720 107692
rect 203760 107652 203766 107664
rect 204714 107652 204720 107664
rect 204772 107652 204778 107704
rect 211798 107652 211804 107704
rect 211856 107692 211862 107704
rect 212810 107692 212816 107704
rect 211856 107664 212816 107692
rect 211856 107652 211862 107664
rect 212810 107652 212816 107664
rect 212868 107652 212874 107704
rect 213178 107652 213184 107704
rect 213236 107692 213242 107704
rect 214098 107692 214104 107704
rect 213236 107664 214104 107692
rect 213236 107652 213242 107664
rect 214098 107652 214104 107664
rect 214156 107652 214162 107704
rect 214650 107652 214656 107704
rect 214708 107692 214714 107704
rect 216122 107692 216128 107704
rect 214708 107664 216128 107692
rect 214708 107652 214714 107664
rect 216122 107652 216128 107664
rect 216180 107652 216186 107704
rect 217318 107652 217324 107704
rect 217376 107692 217382 107704
rect 218146 107692 218152 107704
rect 217376 107664 218152 107692
rect 217376 107652 217382 107664
rect 218146 107652 218152 107664
rect 218204 107652 218210 107704
rect 221550 107652 221556 107704
rect 221608 107692 221614 107704
rect 223022 107692 223028 107704
rect 221608 107664 223028 107692
rect 221608 107652 221614 107664
rect 223022 107652 223028 107664
rect 223080 107652 223086 107704
rect 235442 107652 235448 107704
rect 235500 107692 235506 107704
rect 236362 107692 236368 107704
rect 235500 107664 236368 107692
rect 235500 107652 235506 107664
rect 236362 107652 236368 107664
rect 236420 107652 236426 107704
rect 236638 107652 236644 107704
rect 236696 107692 236702 107704
rect 238386 107692 238392 107704
rect 236696 107664 238392 107692
rect 236696 107652 236702 107664
rect 238386 107652 238392 107664
rect 238444 107652 238450 107704
rect 242158 107652 242164 107704
rect 242216 107692 242222 107704
rect 244918 107692 244924 107704
rect 242216 107664 244924 107692
rect 242216 107652 242222 107664
rect 244918 107652 244924 107664
rect 244976 107652 244982 107704
rect 250530 107652 250536 107704
rect 250588 107692 250594 107704
rect 253382 107692 253388 107704
rect 250588 107664 253388 107692
rect 250588 107652 250594 107664
rect 253382 107652 253388 107664
rect 253440 107652 253446 107704
rect 256050 107652 256056 107704
rect 256108 107692 256114 107704
rect 257062 107692 257068 107704
rect 256108 107664 257068 107692
rect 256108 107652 256114 107664
rect 257062 107652 257068 107664
rect 257120 107652 257126 107704
rect 264238 107652 264244 107704
rect 264296 107692 264302 107704
rect 265158 107692 265164 107704
rect 264296 107664 265164 107692
rect 264296 107652 264302 107664
rect 265158 107652 265164 107664
rect 265216 107652 265222 107704
rect 268378 107652 268384 107704
rect 268436 107692 268442 107704
rect 269206 107692 269212 107704
rect 268436 107664 269212 107692
rect 268436 107652 268442 107664
rect 269206 107652 269212 107664
rect 269264 107652 269270 107704
rect 269758 107652 269764 107704
rect 269816 107692 269822 107704
rect 270494 107692 270500 107704
rect 269816 107664 270500 107692
rect 269816 107652 269822 107664
rect 270494 107652 270500 107664
rect 270552 107652 270558 107704
rect 271138 107652 271144 107704
rect 271196 107692 271202 107704
rect 272058 107692 272064 107704
rect 271196 107664 272064 107692
rect 271196 107652 271202 107664
rect 272058 107652 272064 107664
rect 272116 107652 272122 107704
rect 289078 107652 289084 107704
rect 289136 107692 289142 107704
rect 289906 107692 289912 107704
rect 289136 107664 289912 107692
rect 289136 107652 289142 107664
rect 289906 107652 289912 107664
rect 289964 107652 289970 107704
rect 292390 107652 292396 107704
rect 292448 107692 292454 107704
rect 292666 107692 292672 107704
rect 292448 107664 292672 107692
rect 292448 107652 292454 107664
rect 292666 107652 292672 107664
rect 292724 107652 292730 107704
rect 294782 107652 294788 107704
rect 294840 107692 294846 107704
rect 295978 107692 295984 107704
rect 294840 107664 295984 107692
rect 294840 107652 294846 107664
rect 295978 107652 295984 107664
rect 296036 107652 296042 107704
rect 297266 107652 297272 107704
rect 297324 107692 297330 107704
rect 300026 107692 300032 107704
rect 297324 107664 300032 107692
rect 297324 107652 297330 107664
rect 300026 107652 300032 107664
rect 300084 107652 300090 107704
rect 308214 107652 308220 107704
rect 308272 107692 308278 107704
rect 309962 107692 309968 107704
rect 308272 107664 309968 107692
rect 308272 107652 308278 107664
rect 309962 107652 309968 107664
rect 310020 107652 310026 107704
rect 316678 107652 316684 107704
rect 316736 107692 316742 107704
rect 319438 107692 319444 107704
rect 316736 107664 319444 107692
rect 316736 107652 316742 107664
rect 319438 107652 319444 107664
rect 319496 107652 319502 107704
rect 321554 107652 321560 107704
rect 321612 107692 321618 107704
rect 323578 107692 323584 107704
rect 321612 107664 323584 107692
rect 321612 107652 321618 107664
rect 323578 107652 323584 107664
rect 323636 107652 323642 107704
rect 326430 107652 326436 107704
rect 326488 107692 326494 107704
rect 327810 107692 327816 107704
rect 326488 107664 327816 107692
rect 326488 107652 326494 107664
rect 327810 107652 327816 107664
rect 327868 107652 327874 107704
rect 348326 107652 348332 107704
rect 348384 107692 348390 107704
rect 351178 107692 351184 107704
rect 348384 107664 351184 107692
rect 348384 107652 348390 107664
rect 351178 107652 351184 107664
rect 351236 107652 351242 107704
rect 352006 107652 352012 107704
rect 352064 107692 352070 107704
rect 353938 107692 353944 107704
rect 352064 107664 353944 107692
rect 352064 107652 352070 107664
rect 353938 107652 353944 107664
rect 353996 107652 354002 107704
rect 366634 107652 366640 107704
rect 366692 107692 366698 107704
rect 367738 107692 367744 107704
rect 366692 107664 367744 107692
rect 366692 107652 366698 107664
rect 367738 107652 367744 107664
rect 367796 107652 367802 107704
rect 379974 107652 379980 107704
rect 380032 107692 380038 107704
rect 381538 107692 381544 107704
rect 380032 107664 381544 107692
rect 380032 107652 380038 107664
rect 381538 107652 381544 107664
rect 381596 107652 381602 107704
rect 384022 107652 384028 107704
rect 384080 107692 384086 107704
rect 385678 107692 385684 107704
rect 384080 107664 385684 107692
rect 384080 107652 384086 107664
rect 385678 107652 385684 107664
rect 385736 107652 385742 107704
rect 387334 107652 387340 107704
rect 387392 107692 387398 107704
rect 392670 107692 392676 107704
rect 387392 107664 392676 107692
rect 387392 107652 387398 107664
rect 392670 107652 392676 107664
rect 392728 107652 392734 107704
rect 215386 107108 215392 107160
rect 215444 107148 215450 107160
rect 215570 107148 215576 107160
rect 215444 107120 215576 107148
rect 215444 107108 215450 107120
rect 215570 107108 215576 107120
rect 215628 107108 215634 107160
rect 157334 107040 157340 107092
rect 157392 107080 157398 107092
rect 246114 107080 246120 107092
rect 157392 107052 246120 107080
rect 157392 107040 157398 107052
rect 246114 107040 246120 107052
rect 246172 107040 246178 107092
rect 339862 107040 339868 107092
rect 339920 107080 339926 107092
rect 430574 107080 430580 107092
rect 339920 107052 430580 107080
rect 339920 107040 339926 107052
rect 430574 107040 430580 107052
rect 430632 107040 430638 107092
rect 125594 106972 125600 107024
rect 125652 107012 125658 107024
rect 234890 107012 234896 107024
rect 125652 106984 234896 107012
rect 125652 106972 125658 106984
rect 234890 106972 234896 106984
rect 234948 106972 234954 107024
rect 356882 106972 356888 107024
rect 356940 107012 356946 107024
rect 480254 107012 480260 107024
rect 356940 106984 480260 107012
rect 356940 106972 356946 106984
rect 480254 106972 480260 106984
rect 480312 106972 480318 107024
rect 74534 106904 74540 106956
rect 74592 106944 74598 106956
rect 217686 106944 217692 106956
rect 74592 106916 217692 106944
rect 74592 106904 74598 106916
rect 217686 106904 217692 106916
rect 217744 106904 217750 106956
rect 259454 106904 259460 106956
rect 259512 106944 259518 106956
rect 281442 106944 281448 106956
rect 259512 106916 281448 106944
rect 259512 106904 259518 106916
rect 281442 106904 281448 106916
rect 281500 106904 281506 106956
rect 309410 106904 309416 106956
rect 309468 106944 309474 106956
rect 340874 106944 340880 106956
rect 309468 106916 340880 106944
rect 309468 106904 309474 106916
rect 340874 106904 340880 106916
rect 340932 106904 340938 106956
rect 379606 106904 379612 106956
rect 379664 106944 379670 106956
rect 546494 106944 546500 106956
rect 379664 106916 546500 106944
rect 379664 106904 379670 106916
rect 546494 106904 546500 106916
rect 546552 106904 546558 106956
rect 201494 106836 201500 106888
rect 201552 106876 201558 106888
rect 202046 106876 202052 106888
rect 201552 106848 202052 106876
rect 201552 106836 201558 106848
rect 202046 106836 202052 106848
rect 202104 106836 202110 106888
rect 223758 106836 223764 106888
rect 223816 106876 223822 106888
rect 224310 106876 224316 106888
rect 223816 106848 224316 106876
rect 223816 106836 223822 106848
rect 224310 106836 224316 106848
rect 224368 106836 224374 106888
rect 256878 106836 256884 106888
rect 256936 106876 256942 106888
rect 257614 106876 257620 106888
rect 256936 106848 257620 106876
rect 256936 106836 256942 106848
rect 257614 106836 257620 106848
rect 257672 106836 257678 106888
rect 281718 106836 281724 106888
rect 281776 106876 281782 106888
rect 282270 106876 282276 106888
rect 281776 106848 282276 106876
rect 281776 106836 281782 106848
rect 282270 106836 282276 106848
rect 282328 106836 282334 106888
rect 300854 106836 300860 106888
rect 300912 106876 300918 106888
rect 301406 106876 301412 106888
rect 300912 106848 301412 106876
rect 300912 106836 300918 106848
rect 301406 106836 301412 106848
rect 301464 106836 301470 106888
rect 305086 106836 305092 106888
rect 305144 106876 305150 106888
rect 305822 106876 305828 106888
rect 305144 106848 305828 106876
rect 305144 106836 305150 106848
rect 305822 106836 305828 106848
rect 305880 106836 305886 106888
rect 335354 106836 335360 106888
rect 335412 106876 335418 106888
rect 335906 106876 335912 106888
rect 335412 106848 335912 106876
rect 335412 106836 335418 106848
rect 335906 106836 335912 106848
rect 335964 106836 335970 106888
rect 342254 106836 342260 106888
rect 342312 106876 342318 106888
rect 342806 106876 342812 106888
rect 342312 106848 342812 106876
rect 342312 106836 342318 106848
rect 342806 106836 342812 106848
rect 342864 106836 342870 106888
rect 345106 106836 345112 106888
rect 345164 106876 345170 106888
rect 346026 106876 346032 106888
rect 345164 106848 346032 106876
rect 345164 106836 345170 106848
rect 346026 106836 346032 106848
rect 346084 106836 346090 106888
rect 349338 106836 349344 106888
rect 349396 106876 349402 106888
rect 349614 106876 349620 106888
rect 349396 106848 349620 106876
rect 349396 106836 349402 106848
rect 349614 106836 349620 106848
rect 349672 106836 349678 106888
rect 353386 106836 353392 106888
rect 353444 106876 353450 106888
rect 354122 106876 354128 106888
rect 353444 106848 354128 106876
rect 353444 106836 353450 106848
rect 354122 106836 354128 106848
rect 354180 106836 354186 106888
rect 354766 106836 354772 106888
rect 354824 106876 354830 106888
rect 355318 106876 355324 106888
rect 354824 106848 355324 106876
rect 354824 106836 354830 106848
rect 355318 106836 355324 106848
rect 355376 106836 355382 106888
rect 191834 106768 191840 106820
rect 191892 106808 191898 106820
rect 192662 106808 192668 106820
rect 191892 106780 192668 106808
rect 191892 106768 191898 106780
rect 192662 106768 192668 106780
rect 192720 106768 192726 106820
rect 201586 106768 201592 106820
rect 201644 106808 201650 106820
rect 202414 106808 202420 106820
rect 201644 106780 202420 106808
rect 201644 106768 201650 106780
rect 202414 106768 202420 106780
rect 202472 106768 202478 106820
rect 215386 106768 215392 106820
rect 215444 106808 215450 106820
rect 216214 106808 216220 106820
rect 215444 106780 216220 106808
rect 215444 106768 215450 106780
rect 216214 106768 216220 106780
rect 216272 106768 216278 106820
rect 219434 106768 219440 106820
rect 219492 106808 219498 106820
rect 220262 106808 220268 106820
rect 219492 106780 220268 106808
rect 219492 106768 219498 106780
rect 220262 106768 220268 106780
rect 220320 106768 220326 106820
rect 222286 106768 222292 106820
rect 222344 106808 222350 106820
rect 223114 106808 223120 106820
rect 222344 106780 223120 106808
rect 222344 106768 222350 106780
rect 223114 106768 223120 106780
rect 223172 106768 223178 106820
rect 223666 106768 223672 106820
rect 223724 106808 223730 106820
rect 223942 106808 223948 106820
rect 223724 106780 223948 106808
rect 223724 106768 223730 106780
rect 223942 106768 223948 106780
rect 224000 106768 224006 106820
rect 245746 106768 245752 106820
rect 245804 106808 245810 106820
rect 246574 106808 246580 106820
rect 245804 106780 246580 106808
rect 245804 106768 245810 106780
rect 246574 106768 246580 106780
rect 246632 106768 246638 106820
rect 247126 106768 247132 106820
rect 247184 106808 247190 106820
rect 247862 106808 247868 106820
rect 247184 106780 247868 106808
rect 247184 106768 247190 106780
rect 247862 106768 247868 106780
rect 247920 106768 247926 106820
rect 249886 106768 249892 106820
rect 249944 106808 249950 106820
rect 250714 106808 250720 106820
rect 249944 106780 250720 106808
rect 249944 106768 249950 106780
rect 250714 106768 250720 106780
rect 250772 106768 250778 106820
rect 253934 106768 253940 106820
rect 253992 106808 253998 106820
rect 254762 106808 254768 106820
rect 253992 106780 254768 106808
rect 253992 106768 253998 106780
rect 254762 106768 254768 106780
rect 254820 106768 254826 106820
rect 255314 106768 255320 106820
rect 255372 106808 255378 106820
rect 255958 106808 255964 106820
rect 255372 106780 255964 106808
rect 255372 106768 255378 106780
rect 255958 106768 255964 106780
rect 256016 106768 256022 106820
rect 256786 106768 256792 106820
rect 256844 106808 256850 106820
rect 257154 106808 257160 106820
rect 256844 106780 257160 106808
rect 256844 106768 256850 106780
rect 257154 106768 257160 106780
rect 257212 106768 257218 106820
rect 259546 106768 259552 106820
rect 259604 106808 259610 106820
rect 260374 106808 260380 106820
rect 259604 106780 260380 106808
rect 259604 106768 259610 106780
rect 260374 106768 260380 106780
rect 260432 106768 260438 106820
rect 273346 106768 273352 106820
rect 273404 106808 273410 106820
rect 274174 106808 274180 106820
rect 273404 106780 274180 106808
rect 273404 106768 273410 106780
rect 274174 106768 274180 106780
rect 274232 106768 274238 106820
rect 277578 106768 277584 106820
rect 277636 106808 277642 106820
rect 278222 106808 278228 106820
rect 277636 106780 278228 106808
rect 277636 106768 277642 106780
rect 278222 106768 278228 106780
rect 278280 106768 278286 106820
rect 278866 106768 278872 106820
rect 278924 106808 278930 106820
rect 279510 106808 279516 106820
rect 278924 106780 279516 106808
rect 278924 106768 278930 106780
rect 279510 106768 279516 106780
rect 279568 106768 279574 106820
rect 281626 106768 281632 106820
rect 281684 106808 281690 106820
rect 281902 106808 281908 106820
rect 281684 106780 281908 106808
rect 281684 106768 281690 106780
rect 281902 106768 281908 106780
rect 281960 106768 281966 106820
rect 284386 106768 284392 106820
rect 284444 106808 284450 106820
rect 285214 106808 285220 106820
rect 284444 106780 285220 106808
rect 284444 106768 284450 106780
rect 285214 106768 285220 106780
rect 285272 106768 285278 106820
rect 291194 106768 291200 106820
rect 291252 106808 291258 106820
rect 291654 106808 291660 106820
rect 291252 106780 291660 106808
rect 291252 106768 291258 106780
rect 291654 106768 291660 106780
rect 291712 106768 291718 106820
rect 295426 106768 295432 106820
rect 295484 106808 295490 106820
rect 296070 106808 296076 106820
rect 295484 106780 296076 106808
rect 295484 106768 295490 106780
rect 296070 106768 296076 106780
rect 296128 106768 296134 106820
rect 296806 106768 296812 106820
rect 296864 106808 296870 106820
rect 297726 106808 297732 106820
rect 296864 106780 297732 106808
rect 296864 106768 296870 106780
rect 297726 106768 297732 106780
rect 297784 106768 297790 106820
rect 298094 106768 298100 106820
rect 298152 106808 298158 106820
rect 299014 106808 299020 106820
rect 298152 106780 299020 106808
rect 298152 106768 298158 106780
rect 299014 106768 299020 106780
rect 299072 106768 299078 106820
rect 301038 106768 301044 106820
rect 301096 106808 301102 106820
rect 301774 106808 301780 106820
rect 301096 106780 301780 106808
rect 301096 106768 301102 106780
rect 301774 106768 301780 106780
rect 301832 106768 301838 106820
rect 302234 106768 302240 106820
rect 302292 106808 302298 106820
rect 303062 106808 303068 106820
rect 302292 106780 303068 106808
rect 302292 106768 302298 106780
rect 303062 106768 303068 106780
rect 303120 106768 303126 106820
rect 303706 106768 303712 106820
rect 303764 106808 303770 106820
rect 304258 106808 304264 106820
rect 303764 106780 304264 106808
rect 303764 106768 303770 106780
rect 304258 106768 304264 106780
rect 304316 106768 304322 106820
rect 304994 106768 305000 106820
rect 305052 106808 305058 106820
rect 305454 106808 305460 106820
rect 305052 106780 305460 106808
rect 305052 106768 305058 106780
rect 305454 106768 305460 106780
rect 305512 106768 305518 106820
rect 306374 106768 306380 106820
rect 306432 106808 306438 106820
rect 307110 106808 307116 106820
rect 306432 106780 307116 106808
rect 306432 106768 306438 106780
rect 307110 106768 307116 106780
rect 307168 106768 307174 106820
rect 310514 106768 310520 106820
rect 310572 106808 310578 106820
rect 311526 106808 311532 106820
rect 310572 106780 311532 106808
rect 310572 106768 310578 106780
rect 311526 106768 311532 106780
rect 311584 106768 311590 106820
rect 324314 106768 324320 106820
rect 324372 106808 324378 106820
rect 325326 106808 325332 106820
rect 324372 106780 325332 106808
rect 324372 106768 324378 106780
rect 325326 106768 325332 106780
rect 325384 106768 325390 106820
rect 327166 106768 327172 106820
rect 327224 106808 327230 106820
rect 327718 106808 327724 106820
rect 327224 106780 327724 106808
rect 327224 106768 327230 106780
rect 327718 106768 327724 106780
rect 327776 106768 327782 106820
rect 328546 106768 328552 106820
rect 328604 106808 328610 106820
rect 329374 106808 329380 106820
rect 328604 106780 329380 106808
rect 328604 106768 328610 106780
rect 329374 106768 329380 106780
rect 329432 106768 329438 106820
rect 329834 106768 329840 106820
rect 329892 106808 329898 106820
rect 330662 106808 330668 106820
rect 329892 106780 330668 106808
rect 329892 106768 329898 106780
rect 330662 106768 330668 106780
rect 330720 106768 330726 106820
rect 332594 106768 332600 106820
rect 332652 106808 332658 106820
rect 333422 106808 333428 106820
rect 332652 106780 333428 106808
rect 332652 106768 332658 106780
rect 333422 106768 333428 106780
rect 333480 106768 333486 106820
rect 335538 106768 335544 106820
rect 335596 106808 335602 106820
rect 336274 106808 336280 106820
rect 335596 106780 336280 106808
rect 335596 106768 335602 106780
rect 336274 106768 336280 106780
rect 336332 106768 336338 106820
rect 336734 106768 336740 106820
rect 336792 106808 336798 106820
rect 337102 106808 337108 106820
rect 336792 106780 337108 106808
rect 336792 106768 336798 106780
rect 337102 106768 337108 106780
rect 337160 106768 337166 106820
rect 338206 106768 338212 106820
rect 338264 106808 338270 106820
rect 338758 106808 338764 106820
rect 338264 106780 338764 106808
rect 338264 106768 338270 106780
rect 338758 106768 338764 106780
rect 338816 106768 338822 106820
rect 339494 106768 339500 106820
rect 339552 106808 339558 106820
rect 340322 106808 340328 106820
rect 339552 106780 340328 106808
rect 339552 106768 339558 106780
rect 340322 106768 340328 106780
rect 340380 106768 340386 106820
rect 342438 106768 342444 106820
rect 342496 106808 342502 106820
rect 343174 106808 343180 106820
rect 342496 106780 343180 106808
rect 342496 106768 342502 106780
rect 343174 106768 343180 106780
rect 343232 106768 343238 106820
rect 345198 106768 345204 106820
rect 345256 106808 345262 106820
rect 345566 106808 345572 106820
rect 345256 106780 345572 106808
rect 345256 106768 345262 106780
rect 345566 106768 345572 106780
rect 345624 106768 345630 106820
rect 349154 106768 349160 106820
rect 349212 106808 349218 106820
rect 350074 106808 350080 106820
rect 349212 106780 350080 106808
rect 349212 106768 349218 106780
rect 350074 106768 350080 106780
rect 350132 106768 350138 106820
rect 350534 106768 350540 106820
rect 350592 106808 350598 106820
rect 351270 106808 351276 106820
rect 350592 106780 351276 106808
rect 350592 106768 350598 106780
rect 351270 106768 351276 106780
rect 351328 106768 351334 106820
rect 352006 106768 352012 106820
rect 352064 106808 352070 106820
rect 352926 106808 352932 106820
rect 352064 106780 352932 106808
rect 352064 106768 352070 106780
rect 352926 106768 352932 106780
rect 352984 106768 352990 106820
rect 353294 106768 353300 106820
rect 353352 106808 353358 106820
rect 353754 106808 353760 106820
rect 353352 106780 353760 106808
rect 353352 106768 353358 106780
rect 353754 106768 353760 106780
rect 353812 106768 353818 106820
rect 354674 106768 354680 106820
rect 354732 106808 354738 106820
rect 354950 106808 354956 106820
rect 354732 106780 354956 106808
rect 354732 106768 354738 106780
rect 354950 106768 354956 106780
rect 355008 106768 355014 106820
rect 356054 106768 356060 106820
rect 356112 106808 356118 106820
rect 356238 106808 356244 106820
rect 356112 106780 356244 106808
rect 356112 106768 356118 106780
rect 356238 106768 356244 106780
rect 356296 106768 356302 106820
rect 358814 106768 358820 106820
rect 358872 106808 358878 106820
rect 359826 106808 359832 106820
rect 358872 106780 359832 106808
rect 358872 106768 358878 106780
rect 359826 106768 359832 106780
rect 359884 106768 359890 106820
rect 389266 106768 389272 106820
rect 389324 106808 389330 106820
rect 389818 106808 389824 106820
rect 389324 106780 389824 106808
rect 389324 106768 389330 106780
rect 389818 106768 389824 106780
rect 389876 106768 389882 106820
rect 390554 106768 390560 106820
rect 390612 106808 390618 106820
rect 391474 106808 391480 106820
rect 390612 106780 391480 106808
rect 390612 106768 390618 106780
rect 391474 106768 391480 106780
rect 391532 106768 391538 106820
rect 218238 106700 218244 106752
rect 218296 106740 218302 106752
rect 219066 106740 219072 106752
rect 218296 106712 219072 106740
rect 218296 106700 218302 106712
rect 219066 106700 219072 106712
rect 219124 106700 219130 106752
rect 252738 106700 252744 106752
rect 252796 106740 252802 106752
rect 253566 106740 253572 106752
rect 252796 106712 253572 106740
rect 252796 106700 252802 106712
rect 253566 106700 253572 106712
rect 253624 106700 253630 106752
rect 342346 106700 342352 106752
rect 342404 106740 342410 106752
rect 342622 106740 342628 106752
rect 342404 106712 342628 106740
rect 342404 106700 342410 106712
rect 342622 106700 342628 106712
rect 342680 106700 342686 106752
rect 336826 106632 336832 106684
rect 336884 106672 336890 106684
rect 337470 106672 337476 106684
rect 336884 106644 337476 106672
rect 336884 106632 336890 106644
rect 337470 106632 337476 106644
rect 337528 106632 337534 106684
rect 197446 106088 197452 106140
rect 197504 106128 197510 106140
rect 197998 106128 198004 106140
rect 197504 106100 198004 106128
rect 197504 106088 197510 106100
rect 197998 106088 198004 106100
rect 198056 106088 198062 106140
rect 331214 106088 331220 106140
rect 331272 106128 331278 106140
rect 331398 106128 331404 106140
rect 331272 106100 331404 106128
rect 331272 106088 331278 106100
rect 331398 106088 331404 106100
rect 331456 106088 331462 106140
rect 323026 105816 323032 105868
rect 323084 105856 323090 105868
rect 323670 105856 323676 105868
rect 323084 105828 323676 105856
rect 323084 105816 323090 105828
rect 323670 105816 323676 105828
rect 323728 105816 323734 105868
rect 169754 105680 169760 105732
rect 169812 105720 169818 105732
rect 250622 105720 250628 105732
rect 169812 105692 250628 105720
rect 169812 105680 169818 105692
rect 250622 105680 250628 105692
rect 250680 105680 250686 105732
rect 328914 105680 328920 105732
rect 328972 105720 328978 105732
rect 398834 105720 398840 105732
rect 328972 105692 398840 105720
rect 328972 105680 328978 105692
rect 398834 105680 398840 105692
rect 398892 105680 398898 105732
rect 160094 105612 160100 105664
rect 160152 105652 160158 105664
rect 247310 105652 247316 105664
rect 160152 105624 247316 105652
rect 160152 105612 160158 105624
rect 247310 105612 247316 105624
rect 247368 105612 247374 105664
rect 358078 105612 358084 105664
rect 358136 105652 358142 105664
rect 483014 105652 483020 105664
rect 358136 105624 483020 105652
rect 358136 105612 358142 105624
rect 483014 105612 483020 105624
rect 483072 105612 483078 105664
rect 60734 105544 60740 105596
rect 60792 105584 60798 105596
rect 212902 105584 212908 105596
rect 60792 105556 212908 105584
rect 60792 105544 60798 105556
rect 212902 105544 212908 105556
rect 212960 105544 212966 105596
rect 324406 105544 324412 105596
rect 324464 105584 324470 105596
rect 324590 105584 324596 105596
rect 324464 105556 324596 105584
rect 324464 105544 324470 105556
rect 324590 105544 324596 105556
rect 324648 105544 324654 105596
rect 380434 105544 380440 105596
rect 380492 105584 380498 105596
rect 547874 105584 547880 105596
rect 380492 105556 547880 105584
rect 380492 105544 380498 105556
rect 547874 105544 547880 105556
rect 547932 105544 547938 105596
rect 363230 105408 363236 105460
rect 363288 105448 363294 105460
rect 363506 105448 363512 105460
rect 363288 105420 363512 105448
rect 363288 105408 363294 105420
rect 363506 105408 363512 105420
rect 363564 105408 363570 105460
rect 351914 104728 351920 104780
rect 351972 104768 351978 104780
rect 352558 104768 352564 104780
rect 351972 104740 352564 104768
rect 351972 104728 351978 104740
rect 352558 104728 352564 104740
rect 352616 104728 352622 104780
rect 243078 104592 243084 104644
rect 243136 104592 243142 104644
rect 382366 104592 382372 104644
rect 382424 104592 382430 104644
rect 386598 104592 386604 104644
rect 386656 104592 386662 104644
rect 243096 104440 243124 104592
rect 252554 104456 252560 104508
rect 252612 104496 252618 104508
rect 252830 104496 252836 104508
rect 252612 104468 252836 104496
rect 252612 104456 252618 104468
rect 252830 104456 252836 104468
rect 252888 104456 252894 104508
rect 317506 104456 317512 104508
rect 317564 104496 317570 104508
rect 317690 104496 317696 104508
rect 317564 104468 317696 104496
rect 317564 104456 317570 104468
rect 317690 104456 317696 104468
rect 317748 104456 317754 104508
rect 378134 104456 378140 104508
rect 378192 104496 378198 104508
rect 378410 104496 378416 104508
rect 378192 104468 378416 104496
rect 378192 104456 378198 104468
rect 378410 104456 378416 104468
rect 378468 104456 378474 104508
rect 382384 104440 382412 104592
rect 386616 104440 386644 104592
rect 243078 104388 243084 104440
rect 243136 104388 243142 104440
rect 382366 104388 382372 104440
rect 382424 104388 382430 104440
rect 386598 104388 386604 104440
rect 386656 104388 386662 104440
rect 211430 104320 211436 104372
rect 211488 104360 211494 104372
rect 211614 104360 211620 104372
rect 211488 104332 211620 104360
rect 211488 104320 211494 104332
rect 211614 104320 211620 104332
rect 211672 104320 211678 104372
rect 263870 104320 263876 104372
rect 263928 104360 263934 104372
rect 264054 104360 264060 104372
rect 263928 104332 264060 104360
rect 263928 104320 263934 104332
rect 264054 104320 264060 104332
rect 264112 104320 264118 104372
rect 317414 104320 317420 104372
rect 317472 104360 317478 104372
rect 317598 104360 317604 104372
rect 317472 104332 317604 104360
rect 317472 104320 317478 104332
rect 317598 104320 317604 104332
rect 317656 104320 317662 104372
rect 385126 104320 385132 104372
rect 385184 104360 385190 104372
rect 385770 104360 385776 104372
rect 385184 104332 385776 104360
rect 385184 104320 385190 104332
rect 385770 104320 385776 104332
rect 385828 104320 385834 104372
rect 173894 104252 173900 104304
rect 173952 104292 173958 104304
rect 251818 104292 251824 104304
rect 173952 104264 251824 104292
rect 173952 104252 173958 104264
rect 251818 104252 251824 104264
rect 251876 104252 251882 104304
rect 331306 104252 331312 104304
rect 331364 104292 331370 104304
rect 405734 104292 405740 104304
rect 331364 104264 405740 104292
rect 331364 104252 331370 104264
rect 405734 104252 405740 104264
rect 405792 104252 405798 104304
rect 164234 104184 164240 104236
rect 164292 104224 164298 104236
rect 247218 104224 247224 104236
rect 164292 104196 247224 104224
rect 164292 104184 164298 104196
rect 247218 104184 247224 104196
rect 247276 104184 247282 104236
rect 263686 104184 263692 104236
rect 263744 104224 263750 104236
rect 264422 104224 264428 104236
rect 263744 104196 264428 104224
rect 263744 104184 263750 104196
rect 264422 104184 264428 104196
rect 264480 104184 264486 104236
rect 265066 104184 265072 104236
rect 265124 104224 265130 104236
rect 265710 104224 265716 104236
rect 265124 104196 265716 104224
rect 265124 104184 265130 104196
rect 265710 104184 265716 104196
rect 265768 104184 265774 104236
rect 266538 104184 266544 104236
rect 266596 104224 266602 104236
rect 267366 104224 267372 104236
rect 266596 104196 267372 104224
rect 266596 104184 266602 104196
rect 267366 104184 267372 104196
rect 267424 104184 267430 104236
rect 270678 104184 270684 104236
rect 270736 104224 270742 104236
rect 271414 104224 271420 104236
rect 270736 104196 271420 104224
rect 270736 104184 270742 104196
rect 271414 104184 271420 104196
rect 271472 104184 271478 104236
rect 271966 104184 271972 104236
rect 272024 104224 272030 104236
rect 272610 104224 272616 104236
rect 272024 104196 272616 104224
rect 272024 104184 272030 104196
rect 272610 104184 272616 104196
rect 272668 104184 272674 104236
rect 277394 104184 277400 104236
rect 277452 104224 277458 104236
rect 277854 104224 277860 104236
rect 277452 104196 277860 104224
rect 277452 104184 277458 104196
rect 277854 104184 277860 104196
rect 277912 104184 277918 104236
rect 313366 104184 313372 104236
rect 313424 104224 313430 104236
rect 313918 104224 313924 104236
rect 313424 104196 313924 104224
rect 313424 104184 313430 104196
rect 313918 104184 313924 104196
rect 313976 104184 313982 104236
rect 314654 104184 314660 104236
rect 314712 104224 314718 104236
rect 315206 104224 315212 104236
rect 314712 104196 315212 104224
rect 314712 104184 314718 104196
rect 315206 104184 315212 104196
rect 315264 104184 315270 104236
rect 317414 104184 317420 104236
rect 317472 104224 317478 104236
rect 318058 104224 318064 104236
rect 317472 104196 318064 104224
rect 317472 104184 317478 104196
rect 318058 104184 318064 104196
rect 318116 104184 318122 104236
rect 359274 104184 359280 104236
rect 359332 104224 359338 104236
rect 487154 104224 487160 104236
rect 359332 104196 487160 104224
rect 359332 104184 359338 104196
rect 487154 104184 487160 104196
rect 487212 104184 487218 104236
rect 57974 104116 57980 104168
rect 58032 104156 58038 104168
rect 58032 104128 206968 104156
rect 58032 104116 58038 104128
rect 205634 104048 205640 104100
rect 205692 104088 205698 104100
rect 206462 104088 206468 104100
rect 205692 104060 206468 104088
rect 205692 104048 205698 104060
rect 206462 104048 206468 104060
rect 206520 104048 206526 104100
rect 206940 104088 206968 104128
rect 207014 104116 207020 104168
rect 207072 104156 207078 104168
rect 207658 104156 207664 104168
rect 207072 104128 207664 104156
rect 207072 104116 207078 104128
rect 207658 104116 207664 104128
rect 207716 104116 207722 104168
rect 209774 104116 209780 104168
rect 209832 104156 209838 104168
rect 210510 104156 210516 104168
rect 209832 104128 210516 104156
rect 209832 104116 209838 104128
rect 210510 104116 210516 104128
rect 210568 104116 210574 104168
rect 211246 104116 211252 104168
rect 211304 104156 211310 104168
rect 212166 104156 212172 104168
rect 211304 104128 212172 104156
rect 211304 104116 211310 104128
rect 212166 104116 212172 104128
rect 212224 104116 212230 104168
rect 214006 104116 214012 104168
rect 214064 104156 214070 104168
rect 214558 104156 214564 104168
rect 214064 104128 214564 104156
rect 214064 104116 214070 104128
rect 214558 104116 214564 104128
rect 214616 104116 214622 104168
rect 225046 104116 225052 104168
rect 225104 104156 225110 104168
rect 225598 104156 225604 104168
rect 225104 104128 225604 104156
rect 225104 104116 225110 104128
rect 225598 104116 225604 104128
rect 225656 104116 225662 104168
rect 227714 104116 227720 104168
rect 227772 104156 227778 104168
rect 228358 104156 228364 104168
rect 227772 104128 228364 104156
rect 227772 104116 227778 104128
rect 228358 104116 228364 104128
rect 228416 104116 228422 104168
rect 229278 104116 229284 104168
rect 229336 104156 229342 104168
rect 230014 104156 230020 104168
rect 229336 104128 230020 104156
rect 229336 104116 229342 104128
rect 230014 104116 230020 104128
rect 230072 104116 230078 104168
rect 232038 104116 232044 104168
rect 232096 104156 232102 104168
rect 232406 104156 232412 104168
rect 232096 104128 232412 104156
rect 232096 104116 232102 104128
rect 232406 104116 232412 104128
rect 232464 104116 232470 104168
rect 233326 104116 233332 104168
rect 233384 104156 233390 104168
rect 234062 104156 234068 104168
rect 233384 104128 234068 104156
rect 233384 104116 233390 104128
rect 234062 104116 234068 104128
rect 234120 104116 234126 104168
rect 238846 104116 238852 104168
rect 238904 104156 238910 104168
rect 239306 104156 239312 104168
rect 238904 104128 239312 104156
rect 238904 104116 238910 104128
rect 239306 104116 239312 104128
rect 239364 104116 239370 104168
rect 242986 104116 242992 104168
rect 243044 104156 243050 104168
rect 243814 104156 243820 104168
rect 243044 104128 243820 104156
rect 243044 104116 243050 104128
rect 243814 104116 243820 104128
rect 243872 104116 243878 104168
rect 247034 104116 247040 104168
rect 247092 104156 247098 104168
rect 276934 104156 276940 104168
rect 247092 104128 276940 104156
rect 247092 104116 247098 104128
rect 276934 104116 276940 104128
rect 276992 104116 276998 104168
rect 363046 104116 363052 104168
rect 363104 104156 363110 104168
rect 363414 104156 363420 104168
rect 363104 104128 363420 104156
rect 363104 104116 363110 104128
rect 363414 104116 363420 104128
rect 363472 104116 363478 104168
rect 364334 104116 364340 104168
rect 364392 104156 364398 104168
rect 364702 104156 364708 104168
rect 364392 104128 364708 104156
rect 364392 104116 364398 104128
rect 364702 104116 364708 104128
rect 364760 104116 364766 104168
rect 367094 104116 367100 104168
rect 367152 104156 367158 104168
rect 367554 104156 367560 104168
rect 367152 104128 367560 104156
rect 367152 104116 367158 104128
rect 367554 104116 367560 104128
rect 367612 104116 367618 104168
rect 369854 104116 369860 104168
rect 369912 104156 369918 104168
rect 370774 104156 370780 104168
rect 369912 104128 370780 104156
rect 369912 104116 369918 104128
rect 370774 104116 370780 104128
rect 370832 104116 370838 104168
rect 371234 104116 371240 104168
rect 371292 104156 371298 104168
rect 371970 104156 371976 104168
rect 371292 104128 371976 104156
rect 371292 104116 371298 104128
rect 371970 104116 371976 104128
rect 372028 104116 372034 104168
rect 372614 104116 372620 104168
rect 372672 104156 372678 104168
rect 373626 104156 373632 104168
rect 372672 104128 373632 104156
rect 372672 104116 372678 104128
rect 373626 104116 373632 104128
rect 373684 104116 373690 104168
rect 373994 104116 374000 104168
rect 374052 104156 374058 104168
rect 374822 104156 374828 104168
rect 374052 104128 374828 104156
rect 374052 104116 374058 104128
rect 374822 104116 374828 104128
rect 374880 104116 374886 104168
rect 376754 104116 376760 104168
rect 376812 104156 376818 104168
rect 377214 104156 377220 104168
rect 376812 104128 377220 104156
rect 376812 104116 376818 104128
rect 377214 104116 377220 104128
rect 377272 104116 377278 104168
rect 378226 104116 378232 104168
rect 378284 104156 378290 104168
rect 378870 104156 378876 104168
rect 378284 104128 378876 104156
rect 378284 104116 378290 104128
rect 378870 104116 378876 104128
rect 378928 104116 378934 104168
rect 539594 104156 539600 104168
rect 379486 104128 539600 104156
rect 212074 104088 212080 104100
rect 206940 104060 212080 104088
rect 212074 104048 212080 104060
rect 212132 104048 212138 104100
rect 231946 104048 231952 104100
rect 232004 104088 232010 104100
rect 232774 104088 232780 104100
rect 232004 104060 232780 104088
rect 232004 104048 232010 104060
rect 232774 104048 232780 104060
rect 232832 104048 232838 104100
rect 362954 104048 362960 104100
rect 363012 104088 363018 104100
rect 363874 104088 363880 104100
rect 363012 104060 363880 104088
rect 363012 104048 363018 104060
rect 363874 104048 363880 104060
rect 363932 104048 363938 104100
rect 364426 104048 364432 104100
rect 364484 104088 364490 104100
rect 365070 104088 365076 104100
rect 364484 104060 365076 104088
rect 364484 104048 364490 104060
rect 365070 104048 365076 104060
rect 365128 104048 365134 104100
rect 377122 104048 377128 104100
rect 377180 104088 377186 104100
rect 379486 104088 379514 104128
rect 539594 104116 539600 104128
rect 539652 104116 539658 104168
rect 377180 104060 379514 104088
rect 377180 104048 377186 104060
rect 385034 104048 385040 104100
rect 385092 104088 385098 104100
rect 385402 104088 385408 104100
rect 385092 104060 385408 104088
rect 385092 104048 385098 104060
rect 385402 104048 385408 104060
rect 385460 104048 385466 104100
rect 386506 104048 386512 104100
rect 386564 104088 386570 104100
rect 387426 104088 387432 104100
rect 386564 104060 387432 104088
rect 386564 104048 386570 104060
rect 387426 104048 387432 104060
rect 387484 104048 387490 104100
rect 387978 104048 387984 104100
rect 388036 104088 388042 104100
rect 388622 104088 388628 104100
rect 388036 104060 388628 104088
rect 388036 104048 388042 104060
rect 388622 104048 388628 104060
rect 388680 104048 388686 104100
rect 299474 103912 299480 103964
rect 299532 103952 299538 103964
rect 300118 103952 300124 103964
rect 299532 103924 300124 103952
rect 299532 103912 299538 103924
rect 300118 103912 300124 103924
rect 300176 103912 300182 103964
rect 276014 103504 276020 103556
rect 276072 103544 276078 103556
rect 276198 103544 276204 103556
rect 276072 103516 276204 103544
rect 276072 103504 276078 103516
rect 276198 103504 276204 103516
rect 276256 103504 276262 103556
rect 187694 102892 187700 102944
rect 187752 102932 187758 102944
rect 256970 102932 256976 102944
rect 187752 102904 256976 102932
rect 187752 102892 187758 102904
rect 256970 102892 256976 102904
rect 257028 102892 257034 102944
rect 171134 102824 171140 102876
rect 171192 102864 171198 102876
rect 249886 102864 249892 102876
rect 171192 102836 249892 102864
rect 171192 102824 171198 102836
rect 249886 102824 249892 102836
rect 249944 102824 249950 102876
rect 349430 102824 349436 102876
rect 349488 102864 349494 102876
rect 458174 102864 458180 102876
rect 349488 102836 458180 102864
rect 349488 102824 349494 102836
rect 458174 102824 458180 102836
rect 458232 102824 458238 102876
rect 46934 102756 46940 102808
rect 46992 102796 46998 102808
rect 208302 102796 208308 102808
rect 46992 102768 208308 102796
rect 46992 102756 46998 102768
rect 208302 102756 208308 102768
rect 208360 102756 208366 102808
rect 360286 102756 360292 102808
rect 360344 102796 360350 102808
rect 489914 102796 489920 102808
rect 360344 102768 489920 102796
rect 360344 102756 360350 102768
rect 489914 102756 489920 102768
rect 489972 102756 489978 102808
rect 361574 102144 361580 102196
rect 361632 102184 361638 102196
rect 362310 102184 362316 102196
rect 361632 102156 362316 102184
rect 361632 102144 361638 102156
rect 362310 102144 362316 102156
rect 362368 102144 362374 102196
rect 175274 101532 175280 101584
rect 175332 101572 175338 101584
rect 251358 101572 251364 101584
rect 175332 101544 251364 101572
rect 175332 101532 175338 101544
rect 251358 101532 251364 101544
rect 251416 101532 251422 101584
rect 131114 101464 131120 101516
rect 131172 101504 131178 101516
rect 236914 101504 236920 101516
rect 131172 101476 236920 101504
rect 131172 101464 131178 101476
rect 236914 101464 236920 101476
rect 236972 101464 236978 101516
rect 361758 101464 361764 101516
rect 361816 101504 361822 101516
rect 494054 101504 494060 101516
rect 361816 101476 494060 101504
rect 361816 101464 361822 101476
rect 494054 101464 494060 101476
rect 494112 101464 494118 101516
rect 14458 101396 14464 101448
rect 14516 101436 14522 101448
rect 194686 101436 194692 101448
rect 14516 101408 194692 101436
rect 14516 101396 14522 101408
rect 194686 101396 194692 101408
rect 194744 101396 194750 101448
rect 225138 101396 225144 101448
rect 225196 101436 225202 101448
rect 225966 101436 225972 101448
rect 225196 101408 225972 101436
rect 225196 101396 225202 101408
rect 225966 101396 225972 101408
rect 226024 101396 226030 101448
rect 230382 101396 230388 101448
rect 230440 101436 230446 101448
rect 230566 101436 230572 101448
rect 230440 101408 230572 101436
rect 230440 101396 230446 101408
rect 230566 101396 230572 101408
rect 230624 101396 230630 101448
rect 242894 101396 242900 101448
rect 242952 101436 242958 101448
rect 243170 101436 243176 101448
rect 242952 101408 243176 101436
rect 242952 101396 242958 101408
rect 243170 101396 243176 101408
rect 243228 101396 243234 101448
rect 251174 101396 251180 101448
rect 251232 101436 251238 101448
rect 277394 101436 277400 101448
rect 251232 101408 277400 101436
rect 251232 101396 251238 101408
rect 277394 101396 277400 101408
rect 277452 101396 277458 101448
rect 315574 101396 315580 101448
rect 315632 101436 315638 101448
rect 360286 101436 360292 101448
rect 315632 101408 360292 101436
rect 315632 101396 315638 101408
rect 360286 101396 360292 101408
rect 360344 101396 360350 101448
rect 368474 101396 368480 101448
rect 368532 101436 368538 101448
rect 368658 101436 368664 101448
rect 368532 101408 368664 101436
rect 368532 101396 368538 101408
rect 368658 101396 368664 101408
rect 368716 101396 368722 101448
rect 375466 101396 375472 101448
rect 375524 101436 375530 101448
rect 534074 101436 534080 101448
rect 375524 101408 534080 101436
rect 375524 101396 375530 101408
rect 534074 101396 534080 101408
rect 534132 101396 534138 101448
rect 382274 101328 382280 101380
rect 382332 101368 382338 101380
rect 382458 101368 382464 101380
rect 382332 101340 382464 101368
rect 382332 101328 382338 101340
rect 382458 101328 382464 101340
rect 382516 101328 382522 101380
rect 229186 100920 229192 100972
rect 229244 100960 229250 100972
rect 229462 100960 229468 100972
rect 229244 100932 229468 100960
rect 229244 100920 229250 100932
rect 229462 100920 229468 100932
rect 229520 100920 229526 100972
rect 238938 100716 238944 100768
rect 238996 100756 239002 100768
rect 239766 100756 239772 100768
rect 238996 100728 239772 100756
rect 238996 100716 239002 100728
rect 239766 100716 239772 100728
rect 239824 100716 239830 100768
rect 394418 100648 394424 100700
rect 394476 100688 394482 100700
rect 580166 100688 580172 100700
rect 394476 100660 580172 100688
rect 394476 100648 394482 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 178034 100104 178040 100156
rect 178092 100144 178098 100156
rect 250530 100144 250536 100156
rect 178092 100116 250536 100144
rect 178092 100104 178098 100116
rect 250530 100104 250536 100116
rect 250588 100104 250594 100156
rect 151814 100036 151820 100088
rect 151872 100076 151878 100088
rect 244366 100076 244372 100088
rect 151872 100048 244372 100076
rect 151872 100036 151878 100048
rect 244366 100036 244372 100048
rect 244424 100036 244430 100088
rect 327258 100036 327264 100088
rect 327316 100076 327322 100088
rect 394694 100076 394700 100088
rect 327316 100048 394700 100076
rect 327316 100036 327322 100048
rect 394694 100036 394700 100048
rect 394752 100036 394758 100088
rect 28994 99968 29000 100020
rect 29052 100008 29058 100020
rect 201494 100008 201500 100020
rect 29052 99980 201500 100008
rect 29052 99968 29058 99980
rect 201494 99968 201500 99980
rect 201552 99968 201558 100020
rect 347866 99968 347872 100020
rect 347924 100008 347930 100020
rect 456886 100008 456892 100020
rect 347924 99980 456892 100008
rect 347924 99968 347930 99980
rect 456886 99968 456892 99980
rect 456944 99968 456950 100020
rect 386414 99696 386420 99748
rect 386472 99736 386478 99748
rect 386690 99736 386696 99748
rect 386472 99708 386696 99736
rect 386472 99696 386478 99708
rect 386690 99696 386696 99708
rect 386748 99696 386754 99748
rect 236086 99220 236092 99272
rect 236144 99260 236150 99272
rect 236454 99260 236460 99272
rect 236144 99232 236460 99260
rect 236144 99220 236150 99232
rect 236454 99220 236460 99232
rect 236512 99220 236518 99272
rect 182174 98744 182180 98796
rect 182232 98784 182238 98796
rect 254118 98784 254124 98796
rect 182232 98756 254124 98784
rect 182232 98744 182238 98756
rect 254118 98744 254124 98756
rect 254176 98744 254182 98796
rect 329926 98744 329932 98796
rect 329984 98784 329990 98796
rect 402974 98784 402980 98796
rect 329984 98756 402980 98784
rect 329984 98744 329990 98756
rect 402974 98744 402980 98756
rect 403032 98744 403038 98796
rect 81434 98676 81440 98728
rect 81492 98716 81498 98728
rect 219618 98716 219624 98728
rect 81492 98688 219624 98716
rect 81492 98676 81498 98688
rect 219618 98676 219624 98688
rect 219676 98676 219682 98728
rect 363506 98676 363512 98728
rect 363564 98716 363570 98728
rect 498194 98716 498200 98728
rect 363564 98688 498200 98716
rect 363564 98676 363570 98688
rect 498194 98676 498200 98688
rect 498252 98676 498258 98728
rect 6914 98608 6920 98660
rect 6972 98648 6978 98660
rect 193950 98648 193956 98660
rect 6972 98620 193956 98648
rect 6972 98608 6978 98620
rect 193950 98608 193956 98620
rect 194008 98608 194014 98660
rect 382458 98608 382464 98660
rect 382516 98648 382522 98660
rect 556154 98648 556160 98660
rect 382516 98620 556160 98648
rect 382516 98608 382522 98620
rect 556154 98608 556160 98620
rect 556212 98608 556218 98660
rect 184934 97384 184940 97436
rect 184992 97424 184998 97436
rect 255498 97424 255504 97436
rect 184992 97396 255504 97424
rect 184992 97384 184998 97396
rect 255498 97384 255504 97396
rect 255556 97384 255562 97436
rect 142154 97316 142160 97368
rect 142212 97356 142218 97368
rect 240226 97356 240232 97368
rect 142212 97328 240232 97356
rect 142212 97316 142218 97328
rect 240226 97316 240232 97328
rect 240284 97316 240290 97368
rect 343634 97316 343640 97368
rect 343692 97356 343698 97368
rect 441614 97356 441620 97368
rect 343692 97328 441620 97356
rect 343692 97316 343698 97328
rect 441614 97316 441620 97328
rect 441672 97316 441678 97368
rect 8294 97248 8300 97300
rect 8352 97288 8358 97300
rect 193858 97288 193864 97300
rect 8352 97260 193864 97288
rect 8352 97248 8358 97260
rect 193858 97248 193864 97260
rect 193916 97248 193922 97300
rect 367738 97248 367744 97300
rect 367796 97288 367802 97300
rect 507854 97288 507860 97300
rect 367796 97260 507860 97288
rect 367796 97248 367802 97260
rect 507854 97248 507860 97260
rect 507912 97248 507918 97300
rect 193398 96024 193404 96076
rect 193456 96064 193462 96076
rect 257430 96064 257436 96076
rect 193456 96036 257436 96064
rect 193456 96024 193462 96036
rect 257430 96024 257436 96036
rect 257488 96024 257494 96076
rect 328730 96024 328736 96076
rect 328788 96064 328794 96076
rect 398926 96064 398932 96076
rect 328788 96036 398932 96064
rect 328788 96024 328794 96036
rect 398926 96024 398932 96036
rect 398984 96024 398990 96076
rect 129734 95956 129740 96008
rect 129792 95996 129798 96008
rect 236086 95996 236092 96008
rect 129792 95968 236092 95996
rect 129792 95956 129798 95968
rect 236086 95956 236092 95968
rect 236144 95956 236150 96008
rect 336918 95956 336924 96008
rect 336976 95996 336982 96008
rect 422294 95996 422300 96008
rect 336976 95968 422300 95996
rect 336976 95956 336982 95968
rect 422294 95956 422300 95968
rect 422352 95956 422358 96008
rect 34514 95888 34520 95940
rect 34572 95928 34578 95940
rect 203058 95928 203064 95940
rect 34572 95900 203064 95928
rect 34572 95888 34578 95900
rect 203058 95888 203064 95900
rect 203116 95888 203122 95940
rect 375466 95888 375472 95940
rect 375524 95928 375530 95940
rect 536834 95928 536840 95940
rect 375524 95900 536840 95928
rect 375524 95888 375530 95900
rect 536834 95888 536840 95900
rect 536892 95888 536898 95940
rect 128354 94528 128360 94580
rect 128412 94568 128418 94580
rect 235442 94568 235448 94580
rect 128412 94540 235448 94568
rect 128412 94528 128418 94540
rect 235442 94528 235448 94540
rect 235500 94528 235506 94580
rect 352098 94528 352104 94580
rect 352156 94568 352162 94580
rect 466454 94568 466460 94580
rect 352156 94540 466460 94568
rect 352156 94528 352162 94540
rect 466454 94528 466460 94540
rect 466512 94528 466518 94580
rect 78674 94460 78680 94512
rect 78732 94500 78738 94512
rect 218238 94500 218244 94512
rect 78732 94472 218244 94500
rect 78732 94460 78738 94472
rect 218238 94460 218244 94472
rect 218296 94460 218302 94512
rect 321738 94460 321744 94512
rect 321796 94500 321802 94512
rect 380986 94500 380992 94512
rect 321796 94472 380992 94500
rect 321796 94460 321802 94472
rect 380986 94460 380992 94472
rect 381044 94460 381050 94512
rect 381538 94460 381544 94512
rect 381596 94500 381602 94512
rect 547966 94500 547972 94512
rect 381596 94472 547972 94500
rect 381596 94460 381602 94472
rect 547966 94460 547972 94472
rect 548024 94460 548030 94512
rect 325786 93236 325792 93288
rect 325844 93276 325850 93288
rect 391934 93276 391940 93288
rect 325844 93248 391940 93276
rect 325844 93236 325850 93248
rect 391934 93236 391940 93248
rect 391992 93236 391998 93288
rect 132494 93168 132500 93220
rect 132552 93208 132558 93220
rect 237466 93208 237472 93220
rect 132552 93180 237472 93208
rect 132552 93168 132558 93180
rect 237466 93168 237472 93180
rect 237524 93168 237530 93220
rect 335630 93168 335636 93220
rect 335688 93208 335694 93220
rect 418154 93208 418160 93220
rect 335688 93180 418160 93208
rect 335688 93168 335694 93180
rect 418154 93168 418160 93180
rect 418212 93168 418218 93220
rect 89714 93100 89720 93152
rect 89772 93140 89778 93152
rect 221458 93140 221464 93152
rect 89772 93112 221464 93140
rect 89772 93100 89778 93112
rect 221458 93100 221464 93112
rect 221516 93100 221522 93152
rect 385770 93100 385776 93152
rect 385828 93140 385834 93152
rect 557534 93140 557540 93152
rect 385828 93112 557540 93140
rect 385828 93100 385834 93112
rect 557534 93100 557540 93112
rect 557592 93100 557598 93152
rect 135254 91808 135260 91860
rect 135312 91848 135318 91860
rect 239030 91848 239036 91860
rect 135312 91820 239036 91848
rect 135312 91808 135318 91820
rect 239030 91808 239036 91820
rect 239088 91808 239094 91860
rect 341150 91808 341156 91860
rect 341208 91848 341214 91860
rect 434714 91848 434720 91860
rect 341208 91820 434720 91848
rect 341208 91808 341214 91820
rect 434714 91808 434720 91820
rect 434772 91808 434778 91860
rect 35894 91740 35900 91792
rect 35952 91780 35958 91792
rect 203610 91780 203616 91792
rect 35952 91752 203616 91780
rect 35952 91740 35958 91752
rect 203610 91740 203616 91752
rect 203668 91740 203674 91792
rect 307846 91740 307852 91792
rect 307904 91780 307910 91792
rect 340966 91780 340972 91792
rect 307904 91752 340972 91780
rect 307904 91740 307910 91752
rect 340966 91740 340972 91752
rect 341024 91740 341030 91792
rect 383746 91740 383752 91792
rect 383804 91780 383810 91792
rect 561674 91780 561680 91792
rect 383804 91752 561680 91780
rect 383804 91740 383810 91752
rect 561674 91740 561680 91752
rect 561732 91740 561738 91792
rect 139394 90380 139400 90432
rect 139452 90420 139458 90432
rect 238938 90420 238944 90432
rect 139452 90392 238944 90420
rect 139452 90380 139458 90392
rect 238938 90380 238944 90392
rect 238996 90380 239002 90432
rect 350718 90380 350724 90432
rect 350776 90420 350782 90432
rect 463694 90420 463700 90432
rect 350776 90392 463700 90420
rect 350776 90380 350782 90392
rect 463694 90380 463700 90392
rect 463752 90380 463758 90432
rect 48314 90312 48320 90364
rect 48372 90352 48378 90364
rect 208486 90352 208492 90364
rect 48372 90324 208492 90352
rect 48372 90312 48378 90324
rect 208486 90312 208492 90324
rect 208544 90312 208550 90364
rect 316126 90312 316132 90364
rect 316184 90352 316190 90364
rect 364518 90352 364524 90364
rect 316184 90324 364524 90352
rect 316184 90312 316190 90324
rect 364518 90312 364524 90324
rect 364576 90312 364582 90364
rect 385126 90312 385132 90364
rect 385184 90352 385190 90364
rect 564434 90352 564440 90364
rect 385184 90324 564440 90352
rect 385184 90312 385190 90324
rect 564434 90312 564440 90324
rect 564492 90312 564498 90364
rect 143534 89020 143540 89072
rect 143592 89060 143598 89072
rect 238110 89060 238116 89072
rect 143592 89032 238116 89060
rect 143592 89020 143598 89032
rect 238110 89020 238116 89032
rect 238168 89020 238174 89072
rect 329834 89020 329840 89072
rect 329892 89060 329898 89072
rect 404354 89060 404360 89072
rect 329892 89032 404360 89060
rect 329892 89020 329898 89032
rect 404354 89020 404360 89032
rect 404412 89020 404418 89072
rect 62114 88952 62120 89004
rect 62172 88992 62178 89004
rect 212718 88992 212724 89004
rect 62172 88964 212724 88992
rect 62172 88952 62178 88964
rect 212718 88952 212724 88964
rect 212776 88952 212782 89004
rect 324590 88952 324596 89004
rect 324648 88992 324654 89004
rect 387794 88992 387800 89004
rect 324648 88964 387800 88992
rect 324648 88952 324654 88964
rect 387794 88952 387800 88964
rect 387852 88952 387858 89004
rect 388070 88952 388076 89004
rect 388128 88992 388134 89004
rect 571978 88992 571984 89004
rect 388128 88964 571984 88992
rect 388128 88952 388134 88964
rect 571978 88952 571984 88964
rect 572036 88952 572042 89004
rect 146294 87660 146300 87712
rect 146352 87700 146358 87712
rect 241698 87700 241704 87712
rect 146352 87672 241704 87700
rect 146352 87660 146358 87672
rect 241698 87660 241704 87672
rect 241756 87660 241762 87712
rect 345290 87660 345296 87712
rect 345348 87700 345354 87712
rect 445754 87700 445760 87712
rect 345348 87672 445760 87700
rect 345348 87660 345354 87672
rect 445754 87660 445760 87672
rect 445812 87660 445818 87712
rect 77294 87592 77300 87644
rect 77352 87632 77358 87644
rect 218146 87632 218152 87644
rect 77352 87604 218152 87632
rect 77352 87592 77358 87604
rect 218146 87592 218152 87604
rect 218204 87592 218210 87644
rect 389358 87592 389364 87644
rect 389416 87632 389422 87644
rect 575474 87632 575480 87644
rect 389416 87604 575480 87632
rect 389416 87592 389422 87604
rect 575474 87592 575480 87604
rect 575532 87592 575538 87644
rect 394326 86912 394332 86964
rect 394384 86952 394390 86964
rect 580166 86952 580172 86964
rect 394384 86924 580172 86952
rect 394384 86912 394390 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 150434 86300 150440 86352
rect 150492 86340 150498 86352
rect 243170 86340 243176 86352
rect 150492 86312 243176 86340
rect 150492 86300 150498 86312
rect 243170 86300 243176 86312
rect 243228 86300 243234 86352
rect 114554 86232 114560 86284
rect 114612 86272 114618 86284
rect 230658 86272 230664 86284
rect 114612 86244 230664 86272
rect 114612 86232 114618 86244
rect 230658 86232 230664 86244
rect 230716 86232 230722 86284
rect 327166 86232 327172 86284
rect 327224 86272 327230 86284
rect 396074 86272 396080 86284
rect 327224 86244 396080 86272
rect 327224 86232 327230 86244
rect 396074 86232 396080 86244
rect 396132 86232 396138 86284
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 190086 85524 190092 85536
rect 3384 85496 190092 85524
rect 3384 85484 3390 85496
rect 190086 85484 190092 85496
rect 190144 85484 190150 85536
rect 179414 84872 179420 84924
rect 179472 84912 179478 84924
rect 252738 84912 252744 84924
rect 179472 84884 252744 84912
rect 179472 84872 179478 84884
rect 252738 84872 252744 84884
rect 252796 84872 252802 84924
rect 337378 84872 337384 84924
rect 337436 84912 337442 84924
rect 401594 84912 401600 84924
rect 337436 84884 401600 84912
rect 337436 84872 337442 84884
rect 401594 84872 401600 84884
rect 401652 84872 401658 84924
rect 92474 84804 92480 84856
rect 92532 84844 92538 84856
rect 223850 84844 223856 84856
rect 92532 84816 223856 84844
rect 92532 84804 92538 84816
rect 223850 84804 223856 84816
rect 223908 84804 223914 84856
rect 361666 84804 361672 84856
rect 361724 84844 361730 84856
rect 495434 84844 495440 84856
rect 361724 84816 495440 84844
rect 361724 84804 361730 84816
rect 495434 84804 495440 84816
rect 495492 84804 495498 84856
rect 153194 83512 153200 83564
rect 153252 83552 153258 83564
rect 242158 83552 242164 83564
rect 153252 83524 242164 83552
rect 153252 83512 153258 83524
rect 242158 83512 242164 83524
rect 242216 83512 242222 83564
rect 331398 83512 331404 83564
rect 331456 83552 331462 83564
rect 408494 83552 408500 83564
rect 331456 83524 408500 83552
rect 331456 83512 331462 83524
rect 408494 83512 408500 83524
rect 408552 83512 408558 83564
rect 102134 83444 102140 83496
rect 102192 83484 102198 83496
rect 226426 83484 226432 83496
rect 102192 83456 226432 83484
rect 102192 83444 102198 83456
rect 226426 83444 226432 83456
rect 226484 83444 226490 83496
rect 369118 83444 369124 83496
rect 369176 83484 369182 83496
rect 506474 83484 506480 83496
rect 369176 83456 506480 83484
rect 369176 83444 369182 83456
rect 506474 83444 506480 83456
rect 506532 83444 506538 83496
rect 126974 82152 126980 82204
rect 127032 82192 127038 82204
rect 234706 82192 234712 82204
rect 127032 82164 234712 82192
rect 127032 82152 127038 82164
rect 234706 82152 234712 82164
rect 234764 82152 234770 82204
rect 334158 82152 334164 82204
rect 334216 82192 334222 82204
rect 415394 82192 415400 82204
rect 334216 82164 415400 82192
rect 334216 82152 334222 82164
rect 415394 82152 415400 82164
rect 415452 82152 415458 82204
rect 56594 82084 56600 82136
rect 56652 82124 56658 82136
rect 211338 82124 211344 82136
rect 56652 82096 211344 82124
rect 56652 82084 56658 82096
rect 211338 82084 211344 82096
rect 211396 82084 211402 82136
rect 365806 82084 365812 82136
rect 365864 82124 365870 82136
rect 509234 82124 509240 82136
rect 365864 82096 509240 82124
rect 365864 82084 365870 82096
rect 509234 82084 509240 82096
rect 509292 82084 509298 82136
rect 161474 80724 161480 80776
rect 161532 80764 161538 80776
rect 247218 80764 247224 80776
rect 161532 80736 247224 80764
rect 161532 80724 161538 80736
rect 247218 80724 247224 80736
rect 247276 80724 247282 80776
rect 338298 80724 338304 80776
rect 338356 80764 338362 80776
rect 426434 80764 426440 80776
rect 338356 80736 426440 80764
rect 338356 80724 338362 80736
rect 426434 80724 426440 80736
rect 426492 80724 426498 80776
rect 66254 80656 66260 80708
rect 66312 80696 66318 80708
rect 214006 80696 214012 80708
rect 66312 80668 214012 80696
rect 66312 80656 66318 80668
rect 214006 80656 214012 80668
rect 214064 80656 214070 80708
rect 370038 80656 370044 80708
rect 370096 80696 370102 80708
rect 520274 80696 520280 80708
rect 370096 80668 520280 80696
rect 370096 80656 370102 80668
rect 520274 80656 520280 80668
rect 520332 80656 520338 80708
rect 165614 79364 165620 79416
rect 165672 79404 165678 79416
rect 248506 79404 248512 79416
rect 165672 79376 248512 79404
rect 165672 79364 165678 79376
rect 248506 79364 248512 79376
rect 248564 79364 248570 79416
rect 342530 79364 342536 79416
rect 342588 79404 342594 79416
rect 437474 79404 437480 79416
rect 342588 79376 437480 79404
rect 342588 79364 342594 79376
rect 437474 79364 437480 79376
rect 437532 79364 437538 79416
rect 18598 79296 18604 79348
rect 18656 79336 18662 79348
rect 197538 79336 197544 79348
rect 18656 79308 197544 79336
rect 18656 79296 18662 79308
rect 197538 79296 197544 79308
rect 197596 79296 197602 79348
rect 369946 79296 369952 79348
rect 370004 79336 370010 79348
rect 517514 79336 517520 79348
rect 370004 79308 517520 79336
rect 370004 79296 370010 79308
rect 517514 79296 517520 79308
rect 517572 79296 517578 79348
rect 254118 78140 254124 78192
rect 254176 78180 254182 78192
rect 279050 78180 279056 78192
rect 254176 78152 279056 78180
rect 254176 78140 254182 78152
rect 279050 78140 279056 78152
rect 279108 78140 279114 78192
rect 183554 78004 183560 78056
rect 183612 78044 183618 78056
rect 253934 78044 253940 78056
rect 183612 78016 253940 78044
rect 183612 78004 183618 78016
rect 253934 78004 253940 78016
rect 253992 78004 253998 78056
rect 342438 78004 342444 78056
rect 342496 78044 342502 78056
rect 440326 78044 440332 78056
rect 342496 78016 440332 78044
rect 342496 78004 342502 78016
rect 440326 78004 440332 78016
rect 440384 78004 440390 78056
rect 75914 77936 75920 77988
rect 75972 77976 75978 77988
rect 217318 77976 217324 77988
rect 75972 77948 217324 77976
rect 75972 77936 75978 77948
rect 217318 77936 217324 77948
rect 217376 77936 217382 77988
rect 369854 77936 369860 77988
rect 369912 77976 369918 77988
rect 521654 77976 521660 77988
rect 369912 77948 521660 77976
rect 369912 77936 369918 77948
rect 521654 77936 521660 77948
rect 521712 77936 521718 77988
rect 133874 76576 133880 76628
rect 133932 76616 133938 76628
rect 237558 76616 237564 76628
rect 133932 76588 237564 76616
rect 133932 76576 133938 76588
rect 237558 76576 237564 76588
rect 237616 76576 237622 76628
rect 343726 76576 343732 76628
rect 343784 76616 343790 76628
rect 444374 76616 444380 76628
rect 343784 76588 444380 76616
rect 343784 76576 343790 76588
rect 444374 76576 444380 76588
rect 444432 76576 444438 76628
rect 63494 76508 63500 76560
rect 63552 76548 63558 76560
rect 213178 76548 213184 76560
rect 63552 76520 213184 76548
rect 63552 76508 63558 76520
rect 213178 76508 213184 76520
rect 213236 76508 213242 76560
rect 309226 76508 309232 76560
rect 309284 76548 309290 76560
rect 343634 76548 343640 76560
rect 309284 76520 343640 76548
rect 309284 76508 309290 76520
rect 343634 76508 343640 76520
rect 343692 76508 343698 76560
rect 372890 76508 372896 76560
rect 372948 76548 372954 76560
rect 528554 76548 528560 76560
rect 372948 76520 528560 76548
rect 372948 76508 372954 76520
rect 528554 76508 528560 76520
rect 528612 76508 528618 76560
rect 147674 75216 147680 75268
rect 147732 75256 147738 75268
rect 243078 75256 243084 75268
rect 147732 75228 243084 75256
rect 147732 75216 147738 75228
rect 243078 75216 243084 75228
rect 243136 75216 243142 75268
rect 345198 75216 345204 75268
rect 345256 75256 345262 75268
rect 448514 75256 448520 75268
rect 345256 75228 448520 75256
rect 345256 75216 345262 75228
rect 448514 75216 448520 75228
rect 448572 75216 448578 75268
rect 52454 75148 52460 75200
rect 52512 75188 52518 75200
rect 209958 75188 209964 75200
rect 52512 75160 209964 75188
rect 52512 75148 52518 75160
rect 209958 75148 209964 75160
rect 210016 75148 210022 75200
rect 375374 75148 375380 75200
rect 375432 75188 375438 75200
rect 535454 75188 535460 75200
rect 375432 75160 535460 75188
rect 375432 75148 375438 75160
rect 535454 75148 535460 75160
rect 535512 75148 535518 75200
rect 151906 73856 151912 73908
rect 151964 73896 151970 73908
rect 242986 73896 242992 73908
rect 151964 73868 242992 73896
rect 151964 73856 151970 73868
rect 242986 73856 242992 73868
rect 243044 73856 243050 73908
rect 351178 73856 351184 73908
rect 351236 73896 351242 73908
rect 455414 73896 455420 73908
rect 351236 73868 455420 73896
rect 351236 73856 351242 73868
rect 455414 73856 455420 73868
rect 455472 73856 455478 73908
rect 49694 73788 49700 73840
rect 49752 73828 49758 73840
rect 208578 73828 208584 73840
rect 49752 73800 208584 73828
rect 49752 73788 49758 73800
rect 208578 73788 208584 73800
rect 208636 73788 208642 73840
rect 311986 73788 311992 73840
rect 312044 73828 312050 73840
rect 350718 73828 350724 73840
rect 312044 73800 350724 73828
rect 312044 73788 312050 73800
rect 350718 73788 350724 73800
rect 350776 73788 350782 73840
rect 378318 73788 378324 73840
rect 378376 73828 378382 73840
rect 542354 73828 542360 73840
rect 378376 73800 542360 73828
rect 378376 73788 378382 73800
rect 542354 73788 542360 73800
rect 542412 73788 542418 73840
rect 394234 73108 394240 73160
rect 394292 73148 394298 73160
rect 579982 73148 579988 73160
rect 394292 73120 579988 73148
rect 394292 73108 394298 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 154574 72496 154580 72548
rect 154632 72536 154638 72548
rect 244458 72536 244464 72548
rect 154632 72508 244464 72536
rect 154632 72496 154638 72508
rect 244458 72496 244464 72508
rect 244516 72496 244522 72548
rect 44174 72428 44180 72480
rect 44232 72468 44238 72480
rect 207198 72468 207204 72480
rect 44232 72440 207204 72468
rect 44232 72428 44238 72440
rect 207198 72428 207204 72440
rect 207256 72428 207262 72480
rect 323118 72428 323124 72480
rect 323176 72468 323182 72480
rect 382458 72468 382464 72480
rect 323176 72440 382464 72468
rect 323176 72428 323182 72440
rect 382458 72428 382464 72440
rect 382516 72428 382522 72480
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 189994 71720 190000 71732
rect 3384 71692 190000 71720
rect 3384 71680 3390 71692
rect 189994 71680 190000 71692
rect 190052 71680 190058 71732
rect 353938 71068 353944 71120
rect 353996 71108 354002 71120
rect 465166 71108 465172 71120
rect 353996 71080 465172 71108
rect 353996 71068 354002 71080
rect 465166 71068 465172 71080
rect 465224 71068 465230 71120
rect 185026 71000 185032 71052
rect 185084 71040 185090 71052
rect 255406 71040 255412 71052
rect 185084 71012 255412 71040
rect 185084 71000 185090 71012
rect 255406 71000 255412 71012
rect 255464 71000 255470 71052
rect 379514 71000 379520 71052
rect 379572 71040 379578 71052
rect 549254 71040 549260 71052
rect 379572 71012 549260 71040
rect 379572 71000 379578 71012
rect 549254 71000 549260 71012
rect 549312 71000 549318 71052
rect 162854 69708 162860 69760
rect 162912 69748 162918 69760
rect 247126 69748 247132 69760
rect 162912 69720 247132 69748
rect 162912 69708 162918 69720
rect 247126 69708 247132 69720
rect 247184 69708 247190 69760
rect 352006 69708 352012 69760
rect 352064 69748 352070 69760
rect 469214 69748 469220 69760
rect 352064 69720 469220 69748
rect 352064 69708 352070 69720
rect 469214 69708 469220 69720
rect 469272 69708 469278 69760
rect 41414 69640 41420 69692
rect 41472 69680 41478 69692
rect 205818 69680 205824 69692
rect 41472 69652 205824 69680
rect 41472 69640 41478 69652
rect 205818 69640 205824 69652
rect 205876 69640 205882 69692
rect 381078 69640 381084 69692
rect 381136 69680 381142 69692
rect 553394 69680 553400 69692
rect 381136 69652 553400 69680
rect 381136 69640 381142 69652
rect 553394 69640 553400 69652
rect 553452 69640 553458 69692
rect 166994 68348 167000 68400
rect 167052 68388 167058 68400
rect 248598 68388 248604 68400
rect 167052 68360 248604 68388
rect 167052 68348 167058 68360
rect 248598 68348 248604 68360
rect 248656 68348 248662 68400
rect 356238 68348 356244 68400
rect 356296 68388 356302 68400
rect 481634 68388 481640 68400
rect 356296 68360 481640 68388
rect 356296 68348 356302 68360
rect 481634 68348 481640 68360
rect 481692 68348 481698 68400
rect 27614 68280 27620 68332
rect 27672 68320 27678 68332
rect 201678 68320 201684 68332
rect 27672 68292 201684 68320
rect 27672 68280 27678 68292
rect 201678 68280 201684 68292
rect 201736 68280 201742 68332
rect 383654 68280 383660 68332
rect 383712 68320 383718 68332
rect 560294 68320 560300 68332
rect 383712 68292 560300 68320
rect 383712 68280 383718 68292
rect 560294 68280 560300 68292
rect 560352 68280 560358 68332
rect 180794 66920 180800 66972
rect 180852 66960 180858 66972
rect 254026 66960 254032 66972
rect 180852 66932 254032 66960
rect 180852 66920 180858 66932
rect 254026 66920 254032 66932
rect 254084 66920 254090 66972
rect 91094 66852 91100 66904
rect 91152 66892 91158 66904
rect 222286 66892 222292 66904
rect 91152 66864 222292 66892
rect 91152 66852 91158 66864
rect 222286 66852 222292 66864
rect 222344 66852 222350 66904
rect 314838 66852 314844 66904
rect 314896 66892 314902 66904
rect 357434 66892 357440 66904
rect 314896 66864 357440 66892
rect 314896 66852 314902 66864
rect 357434 66852 357440 66864
rect 357492 66852 357498 66904
rect 357618 66852 357624 66904
rect 357676 66892 357682 66904
rect 484394 66892 484400 66904
rect 357676 66864 484400 66892
rect 357676 66852 357682 66864
rect 484394 66852 484400 66864
rect 484452 66852 484458 66904
rect 135346 65560 135352 65612
rect 135404 65600 135410 65612
rect 236638 65600 236644 65612
rect 135404 65572 236644 65600
rect 135404 65560 135410 65572
rect 236638 65560 236644 65572
rect 236696 65560 236702 65612
rect 95234 65492 95240 65544
rect 95292 65532 95298 65544
rect 225230 65532 225236 65544
rect 95292 65504 225236 65532
rect 95292 65492 95298 65504
rect 225230 65492 225236 65504
rect 225288 65492 225294 65544
rect 358998 65492 359004 65544
rect 359056 65532 359062 65544
rect 488534 65532 488540 65544
rect 359056 65504 488540 65532
rect 359056 65492 359062 65504
rect 488534 65492 488540 65504
rect 488592 65492 488598 65544
rect 138014 64200 138020 64252
rect 138072 64240 138078 64252
rect 238846 64240 238852 64252
rect 138072 64212 238852 64240
rect 138072 64200 138078 64212
rect 238846 64200 238852 64212
rect 238904 64200 238910 64252
rect 99374 64132 99380 64184
rect 99432 64172 99438 64184
rect 225138 64172 225144 64184
rect 99432 64144 225144 64172
rect 99432 64132 99438 64144
rect 225138 64132 225144 64144
rect 225196 64132 225202 64184
rect 363138 64132 363144 64184
rect 363196 64172 363202 64184
rect 498286 64172 498292 64184
rect 363196 64144 498292 64172
rect 363196 64132 363202 64144
rect 498286 64132 498292 64144
rect 498344 64132 498350 64184
rect 155954 62840 155960 62892
rect 156012 62880 156018 62892
rect 245838 62880 245844 62892
rect 156012 62852 245844 62880
rect 156012 62840 156018 62852
rect 245838 62840 245844 62852
rect 245896 62840 245902 62892
rect 331306 62840 331312 62892
rect 331364 62880 331370 62892
rect 407114 62880 407120 62892
rect 331364 62852 407120 62880
rect 331364 62840 331370 62852
rect 407114 62840 407120 62852
rect 407172 62840 407178 62892
rect 21358 62772 21364 62824
rect 21416 62812 21422 62824
rect 196158 62812 196164 62824
rect 21416 62784 196164 62812
rect 21416 62772 21422 62784
rect 196158 62772 196164 62784
rect 196216 62772 196222 62824
rect 364610 62772 364616 62824
rect 364668 62812 364674 62824
rect 502334 62812 502340 62824
rect 364668 62784 502340 62812
rect 364668 62772 364674 62784
rect 502334 62772 502340 62784
rect 502392 62772 502398 62824
rect 69014 61344 69020 61396
rect 69072 61384 69078 61396
rect 215478 61384 215484 61396
rect 69072 61356 215484 61384
rect 69072 61344 69078 61356
rect 215478 61344 215484 61356
rect 215536 61344 215542 61396
rect 310698 61344 310704 61396
rect 310756 61384 310762 61396
rect 347866 61384 347872 61396
rect 310756 61356 347872 61384
rect 310756 61344 310762 61356
rect 347866 61344 347872 61356
rect 347924 61344 347930 61396
rect 367278 61344 367284 61396
rect 367336 61384 367342 61396
rect 513374 61384 513380 61396
rect 367336 61356 513380 61384
rect 367336 61344 367342 61356
rect 513374 61344 513380 61356
rect 513432 61344 513438 61396
rect 394142 60664 394148 60716
rect 394200 60704 394206 60716
rect 580166 60704 580172 60716
rect 394200 60676 580172 60704
rect 394200 60664 394206 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 71774 59984 71780 60036
rect 71832 60024 71838 60036
rect 216766 60024 216772 60036
rect 71832 59996 216772 60024
rect 71832 59984 71838 59996
rect 216766 59984 216772 59996
rect 216824 59984 216830 60036
rect 328638 59984 328644 60036
rect 328696 60024 328702 60036
rect 397454 60024 397460 60036
rect 328696 59996 397460 60024
rect 328696 59984 328702 59996
rect 397454 59984 397460 59996
rect 397512 59984 397518 60036
rect 85574 58624 85580 58676
rect 85632 58664 85638 58676
rect 220998 58664 221004 58676
rect 85632 58636 221004 58664
rect 85632 58624 85638 58636
rect 220998 58624 221004 58636
rect 221056 58624 221062 58676
rect 317690 58624 317696 58676
rect 317748 58664 317754 58676
rect 368658 58664 368664 58676
rect 317748 58636 368664 58664
rect 317748 58624 317754 58636
rect 368658 58624 368664 58636
rect 368716 58624 368722 58676
rect 368750 58624 368756 58676
rect 368808 58664 368814 58676
rect 516134 58664 516140 58676
rect 368808 58636 516140 58664
rect 368808 58624 368814 58636
rect 516134 58624 516140 58636
rect 516192 58624 516198 58676
rect 328546 57264 328552 57316
rect 328604 57304 328610 57316
rect 400214 57304 400220 57316
rect 328604 57276 400220 57304
rect 328604 57264 328610 57276
rect 400214 57264 400220 57276
rect 400272 57264 400278 57316
rect 100754 57196 100760 57248
rect 100812 57236 100818 57248
rect 220078 57236 220084 57248
rect 100812 57208 220084 57236
rect 100812 57196 100818 57208
rect 220078 57196 220084 57208
rect 220136 57196 220142 57248
rect 385678 57196 385684 57248
rect 385736 57236 385742 57248
rect 558914 57236 558920 57248
rect 385736 57208 558920 57236
rect 385736 57196 385742 57208
rect 558914 57196 558920 57208
rect 558972 57196 558978 57248
rect 110506 55836 110512 55888
rect 110564 55876 110570 55888
rect 229278 55876 229284 55888
rect 110564 55848 229284 55876
rect 110564 55836 110570 55848
rect 229278 55836 229284 55848
rect 229336 55836 229342 55888
rect 324498 55836 324504 55888
rect 324556 55876 324562 55888
rect 385126 55876 385132 55888
rect 324556 55848 385132 55876
rect 324556 55836 324562 55848
rect 385126 55836 385132 55848
rect 385184 55836 385190 55888
rect 385218 55836 385224 55888
rect 385276 55876 385282 55888
rect 563054 55876 563060 55888
rect 385276 55848 563060 55876
rect 385276 55836 385282 55848
rect 563054 55836 563060 55848
rect 563112 55836 563118 55888
rect 160186 54544 160192 54596
rect 160244 54584 160250 54596
rect 245746 54584 245752 54596
rect 160244 54556 245752 54584
rect 160244 54544 160250 54556
rect 245746 54544 245752 54556
rect 245804 54544 245810 54596
rect 324406 54544 324412 54596
rect 324464 54584 324470 54596
rect 386690 54584 386696 54596
rect 324464 54556 386696 54584
rect 324464 54544 324470 54556
rect 386690 54544 386696 54556
rect 386748 54544 386754 54596
rect 88334 54476 88340 54528
rect 88392 54516 88398 54528
rect 222378 54516 222384 54528
rect 88392 54488 222384 54516
rect 88392 54476 88398 54488
rect 222378 54476 222384 54488
rect 222436 54476 222442 54528
rect 386598 54476 386604 54528
rect 386656 54516 386662 54528
rect 565814 54516 565820 54528
rect 386656 54488 565820 54516
rect 386656 54476 386662 54488
rect 565814 54476 565820 54488
rect 565872 54476 565878 54528
rect 149054 53116 149060 53168
rect 149112 53156 149118 53168
rect 242894 53156 242900 53168
rect 149112 53128 242900 53156
rect 149112 53116 149118 53128
rect 242894 53116 242900 53128
rect 242952 53116 242958 53168
rect 102226 53048 102232 53100
rect 102284 53088 102290 53100
rect 226518 53088 226524 53100
rect 102284 53060 226524 53088
rect 102284 53048 102290 53060
rect 226518 53048 226524 53060
rect 226576 53048 226582 53100
rect 321646 53048 321652 53100
rect 321704 53088 321710 53100
rect 379514 53088 379520 53100
rect 321704 53060 379520 53088
rect 321704 53048 321710 53060
rect 379514 53048 379520 53060
rect 379572 53048 379578 53100
rect 386506 53048 386512 53100
rect 386564 53088 386570 53100
rect 569954 53088 569960 53100
rect 386564 53060 569960 53088
rect 386564 53048 386570 53060
rect 569954 53048 569960 53060
rect 570012 53048 570018 53100
rect 219618 51756 219624 51808
rect 219676 51796 219682 51808
rect 266538 51796 266544 51808
rect 219676 51768 266544 51796
rect 219676 51756 219682 51768
rect 266538 51756 266544 51768
rect 266596 51756 266602 51808
rect 121454 51688 121460 51740
rect 121512 51728 121518 51740
rect 233418 51728 233424 51740
rect 121512 51700 233424 51728
rect 121512 51688 121518 51700
rect 233418 51688 233424 51700
rect 233476 51688 233482 51740
rect 320358 51688 320364 51740
rect 320416 51728 320422 51740
rect 375374 51728 375380 51740
rect 320416 51700 375380 51728
rect 320416 51688 320422 51700
rect 375374 51688 375380 51700
rect 375432 51688 375438 51740
rect 387978 51688 387984 51740
rect 388036 51728 388042 51740
rect 572070 51728 572076 51740
rect 388036 51700 572076 51728
rect 388036 51688 388042 51700
rect 572070 51688 572076 51700
rect 572128 51688 572134 51740
rect 144914 50328 144920 50380
rect 144972 50368 144978 50380
rect 241606 50368 241612 50380
rect 144972 50340 241612 50368
rect 144972 50328 144978 50340
rect 241606 50328 241612 50340
rect 241664 50328 241670 50380
rect 317598 50328 317604 50380
rect 317656 50368 317662 50380
rect 365806 50368 365812 50380
rect 317656 50340 365812 50368
rect 317656 50328 317662 50340
rect 365806 50328 365812 50340
rect 365864 50328 365870 50380
rect 389266 50328 389272 50380
rect 389324 50368 389330 50380
rect 574738 50368 574744 50380
rect 389324 50340 574744 50368
rect 389324 50328 389330 50340
rect 574738 50328 574744 50340
rect 574796 50328 574802 50380
rect 346486 49036 346492 49088
rect 346544 49076 346550 49088
rect 452654 49076 452660 49088
rect 346544 49048 452660 49076
rect 346544 49036 346550 49048
rect 452654 49036 452660 49048
rect 452712 49036 452718 49088
rect 59354 48968 59360 49020
rect 59412 49008 59418 49020
rect 211246 49008 211252 49020
rect 59412 48980 211252 49008
rect 59412 48968 59418 48980
rect 211246 48968 211252 48980
rect 211304 48968 211310 49020
rect 216766 48968 216772 49020
rect 216824 49008 216830 49020
rect 266446 49008 266452 49020
rect 216824 48980 266452 49008
rect 216824 48968 216830 48980
rect 266446 48968 266452 48980
rect 266504 48968 266510 49020
rect 389174 48968 389180 49020
rect 389232 49008 389238 49020
rect 574094 49008 574100 49020
rect 389232 48980 574100 49008
rect 389232 48968 389238 48980
rect 574094 48968 574100 48980
rect 574152 48968 574158 49020
rect 209958 47608 209964 47660
rect 210016 47648 210022 47660
rect 263778 47648 263784 47660
rect 210016 47620 263784 47648
rect 210016 47608 210022 47620
rect 263778 47608 263784 47620
rect 263836 47608 263842 47660
rect 349338 47608 349344 47660
rect 349396 47648 349402 47660
rect 459554 47648 459560 47660
rect 349396 47620 459560 47648
rect 349396 47608 349402 47620
rect 459554 47608 459560 47620
rect 459612 47608 459618 47660
rect 86954 47540 86960 47592
rect 87012 47580 87018 47592
rect 218698 47580 218704 47592
rect 87012 47552 218704 47580
rect 87012 47540 87018 47552
rect 218698 47540 218704 47552
rect 218756 47540 218762 47592
rect 400858 47540 400864 47592
rect 400916 47580 400922 47592
rect 578234 47580 578240 47592
rect 400916 47552 578240 47580
rect 400916 47540 400922 47552
rect 578234 47540 578240 47552
rect 578292 47540 578298 47592
rect 143626 46180 143632 46232
rect 143684 46220 143690 46232
rect 241514 46220 241520 46232
rect 143684 46192 241520 46220
rect 143684 46180 143690 46192
rect 241514 46180 241520 46192
rect 241572 46180 241578 46232
rect 353478 46180 353484 46232
rect 353536 46220 353542 46232
rect 470594 46220 470600 46232
rect 353536 46192 470600 46220
rect 353536 46180 353542 46192
rect 470594 46180 470600 46192
rect 470652 46180 470658 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 189902 45540 189908 45552
rect 3568 45512 189908 45540
rect 3568 45500 3574 45512
rect 189902 45500 189908 45512
rect 189960 45500 189966 45552
rect 205818 44820 205824 44872
rect 205876 44860 205882 44872
rect 262306 44860 262312 44872
rect 205876 44832 262312 44860
rect 205876 44820 205882 44832
rect 262306 44820 262312 44832
rect 262364 44820 262370 44872
rect 356146 44820 356152 44872
rect 356204 44860 356210 44872
rect 477494 44860 477500 44872
rect 356204 44832 477500 44860
rect 356204 44820 356210 44832
rect 477494 44820 477500 44832
rect 477552 44820 477558 44872
rect 199010 43460 199016 43512
rect 199068 43500 199074 43512
rect 259730 43500 259736 43512
rect 199068 43472 259736 43500
rect 199068 43460 199074 43472
rect 259730 43460 259736 43472
rect 259788 43460 259794 43512
rect 30374 43392 30380 43444
rect 30432 43432 30438 43444
rect 201586 43432 201592 43444
rect 30432 43404 201592 43432
rect 30432 43392 30438 43404
rect 201586 43392 201592 43404
rect 201644 43392 201650 43444
rect 357526 43392 357532 43444
rect 357584 43432 357590 43444
rect 481726 43432 481732 43444
rect 357584 43404 481732 43432
rect 357584 43392 357590 43404
rect 481726 43392 481732 43404
rect 481784 43392 481790 43444
rect 176654 42100 176660 42152
rect 176712 42140 176718 42152
rect 252646 42140 252652 42152
rect 176712 42112 252652 42140
rect 176712 42100 176718 42112
rect 252646 42100 252652 42112
rect 252704 42100 252710 42152
rect 70394 42032 70400 42084
rect 70452 42072 70458 42084
rect 215386 42072 215392 42084
rect 70452 42044 215392 42072
rect 70452 42032 70458 42044
rect 215386 42032 215392 42044
rect 215444 42032 215450 42084
rect 358906 42032 358912 42084
rect 358964 42072 358970 42084
rect 485774 42072 485780 42084
rect 358964 42044 485780 42072
rect 358964 42032 358970 42044
rect 485774 42032 485780 42044
rect 485832 42032 485838 42084
rect 158714 40672 158720 40724
rect 158772 40712 158778 40724
rect 245930 40712 245936 40724
rect 158772 40684 245936 40712
rect 158772 40672 158778 40684
rect 245930 40672 245936 40684
rect 245988 40672 245994 40724
rect 363046 40672 363052 40724
rect 363104 40712 363110 40724
rect 499574 40712 499580 40724
rect 363104 40684 499580 40712
rect 363104 40672 363110 40684
rect 499574 40672 499580 40684
rect 499632 40672 499638 40724
rect 127066 39312 127072 39364
rect 127124 39352 127130 39364
rect 236270 39352 236276 39364
rect 127124 39324 236276 39352
rect 127124 39312 127130 39324
rect 236270 39312 236276 39324
rect 236328 39312 236334 39364
rect 242894 39312 242900 39364
rect 242952 39352 242958 39364
rect 274910 39352 274916 39364
rect 242952 39324 274916 39352
rect 242952 39312 242958 39324
rect 274910 39312 274916 39324
rect 274968 39312 274974 39364
rect 365714 39312 365720 39364
rect 365772 39352 365778 39364
rect 506566 39352 506572 39364
rect 365772 39324 506572 39352
rect 365772 39312 365778 39324
rect 506566 39312 506572 39324
rect 506624 39312 506630 39364
rect 136634 37884 136640 37936
rect 136692 37924 136698 37936
rect 238754 37924 238760 37936
rect 136692 37896 238760 37924
rect 136692 37884 136698 37896
rect 238754 37884 238760 37896
rect 238812 37884 238818 37936
rect 316034 37884 316040 37936
rect 316092 37924 316098 37936
rect 361666 37924 361672 37936
rect 316092 37896 361672 37924
rect 316092 37884 316098 37896
rect 361666 37884 361672 37896
rect 361724 37884 361730 37936
rect 368566 37884 368572 37936
rect 368624 37924 368630 37936
rect 514754 37924 514760 37936
rect 368624 37896 514760 37924
rect 368624 37884 368630 37896
rect 514754 37884 514760 37896
rect 514812 37884 514818 37936
rect 235994 36592 236000 36644
rect 236052 36632 236058 36644
rect 273438 36632 273444 36644
rect 236052 36604 273444 36632
rect 236052 36592 236058 36604
rect 273438 36592 273444 36604
rect 273496 36592 273502 36644
rect 140774 36524 140780 36576
rect 140832 36564 140838 36576
rect 238018 36564 238024 36576
rect 140832 36536 238024 36564
rect 140832 36524 140838 36536
rect 238018 36524 238024 36536
rect 238076 36524 238082 36576
rect 314746 36524 314752 36576
rect 314804 36564 314810 36576
rect 357526 36564 357532 36576
rect 314804 36536 357532 36564
rect 314804 36524 314810 36536
rect 357526 36524 357532 36536
rect 357584 36524 357590 36576
rect 361574 36524 361580 36576
rect 361632 36564 361638 36576
rect 496814 36564 496820 36576
rect 361632 36536 496820 36564
rect 361632 36524 361638 36536
rect 496814 36524 496820 36536
rect 496872 36524 496878 36576
rect 118694 35164 118700 35216
rect 118752 35204 118758 35216
rect 232038 35204 232044 35216
rect 118752 35176 232044 35204
rect 118752 35164 118758 35176
rect 232038 35164 232044 35176
rect 232096 35164 232102 35216
rect 233418 35164 233424 35216
rect 233476 35204 233482 35216
rect 271138 35204 271144 35216
rect 233476 35176 271144 35204
rect 233476 35164 233482 35176
rect 271138 35164 271144 35176
rect 271196 35164 271202 35216
rect 313458 35164 313464 35216
rect 313516 35204 313522 35216
rect 354950 35204 354956 35216
rect 313516 35176 354956 35204
rect 313516 35164 313522 35176
rect 354950 35164 354956 35176
rect 355008 35164 355014 35216
rect 358814 35164 358820 35216
rect 358872 35204 358878 35216
rect 490006 35204 490012 35216
rect 358872 35176 490012 35204
rect 358872 35164 358878 35176
rect 490006 35164 490012 35176
rect 490064 35164 490070 35216
rect 345106 33804 345112 33856
rect 345164 33844 345170 33856
rect 448606 33844 448612 33856
rect 345164 33816 448612 33844
rect 345164 33804 345170 33816
rect 448606 33804 448612 33816
rect 448664 33804 448670 33856
rect 17954 33736 17960 33788
rect 18012 33776 18018 33788
rect 197446 33776 197452 33788
rect 18012 33748 197452 33776
rect 18012 33736 18018 33748
rect 197446 33736 197452 33748
rect 197504 33736 197510 33788
rect 197538 33736 197544 33788
rect 197596 33776 197602 33788
rect 259638 33776 259644 33788
rect 197596 33748 259644 33776
rect 197596 33736 197602 33748
rect 259638 33736 259644 33748
rect 259696 33736 259702 33788
rect 386414 33736 386420 33788
rect 386472 33776 386478 33788
rect 567194 33776 567200 33788
rect 386472 33748 567200 33776
rect 386472 33736 386478 33748
rect 567194 33736 567200 33748
rect 567252 33736 567258 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 189810 33096 189816 33108
rect 2924 33068 189816 33096
rect 2924 33056 2930 33068
rect 189810 33056 189816 33068
rect 189868 33056 189874 33108
rect 394050 33056 394056 33108
rect 394108 33096 394114 33108
rect 580166 33096 580172 33108
rect 394108 33068 580172 33096
rect 394108 33056 394114 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 189074 32376 189080 32428
rect 189132 32416 189138 32428
rect 255958 32416 255964 32428
rect 189132 32388 255964 32416
rect 189132 32376 189138 32388
rect 255958 32376 255964 32388
rect 256016 32376 256022 32428
rect 324314 32376 324320 32428
rect 324372 32416 324378 32428
rect 389174 32416 389180 32428
rect 324372 32388 389180 32416
rect 324372 32376 324378 32388
rect 389174 32376 389180 32388
rect 389232 32376 389238 32428
rect 215386 31084 215392 31136
rect 215444 31124 215450 31136
rect 265066 31124 265072 31136
rect 215444 31096 265072 31124
rect 215444 31084 215450 31096
rect 265066 31084 265072 31096
rect 265124 31084 265130 31136
rect 73154 31016 73160 31068
rect 73212 31056 73218 31068
rect 216858 31056 216864 31068
rect 73212 31028 216864 31056
rect 73212 31016 73218 31028
rect 216858 31016 216864 31028
rect 216916 31016 216922 31068
rect 307754 31016 307760 31068
rect 307812 31056 307818 31068
rect 336918 31056 336924 31068
rect 307812 31028 336924 31056
rect 307812 31016 307818 31028
rect 336918 31016 336924 31028
rect 336976 31016 336982 31068
rect 371418 31016 371424 31068
rect 371476 31056 371482 31068
rect 523034 31056 523040 31068
rect 371476 31028 523040 31056
rect 371476 31016 371482 31028
rect 523034 31016 523040 31028
rect 523092 31016 523098 31068
rect 193490 29656 193496 29708
rect 193548 29696 193554 29708
rect 258166 29696 258172 29708
rect 193548 29668 258172 29696
rect 193548 29656 193554 29668
rect 258166 29656 258172 29668
rect 258224 29656 258230 29708
rect 338758 29656 338764 29708
rect 338816 29696 338822 29708
rect 411254 29696 411260 29708
rect 338816 29668 411260 29696
rect 338816 29656 338822 29668
rect 411254 29656 411260 29668
rect 411312 29656 411318 29708
rect 60826 29588 60832 29640
rect 60884 29628 60890 29640
rect 211798 29628 211804 29640
rect 60884 29600 211804 29628
rect 60884 29588 60890 29600
rect 211798 29588 211804 29600
rect 211856 29588 211862 29640
rect 311894 29588 311900 29640
rect 311952 29628 311958 29640
rect 349338 29628 349344 29640
rect 311952 29600 349344 29628
rect 311952 29588 311958 29600
rect 349338 29588 349344 29600
rect 349396 29588 349402 29640
rect 395338 29588 395344 29640
rect 395396 29628 395402 29640
rect 580258 29628 580264 29640
rect 395396 29600 580264 29628
rect 395396 29588 395402 29600
rect 580258 29588 580264 29600
rect 580316 29588 580322 29640
rect 310606 28432 310612 28484
rect 310664 28472 310670 28484
rect 346486 28472 346492 28484
rect 310664 28444 346492 28472
rect 310664 28432 310670 28444
rect 346486 28432 346492 28444
rect 346544 28432 346550 28484
rect 190454 28296 190460 28348
rect 190512 28336 190518 28348
rect 256786 28336 256792 28348
rect 190512 28308 256792 28336
rect 190512 28296 190518 28308
rect 256786 28296 256792 28308
rect 256844 28296 256850 28348
rect 346394 28296 346400 28348
rect 346452 28336 346458 28348
rect 451274 28336 451280 28348
rect 346452 28308 451280 28336
rect 346452 28296 346458 28308
rect 451274 28296 451280 28308
rect 451332 28296 451338 28348
rect 67634 28228 67640 28280
rect 67692 28268 67698 28280
rect 215570 28268 215576 28280
rect 67692 28240 215576 28268
rect 67692 28228 67698 28240
rect 215570 28228 215576 28240
rect 215628 28228 215634 28280
rect 387886 28228 387892 28280
rect 387944 28268 387950 28280
rect 570598 28268 570604 28280
rect 387944 28240 570604 28268
rect 387944 28228 387950 28240
rect 570598 28228 570604 28240
rect 570656 28228 570662 28280
rect 186314 26936 186320 26988
rect 186372 26976 186378 26988
rect 255314 26976 255320 26988
rect 186372 26948 255320 26976
rect 186372 26936 186378 26948
rect 255314 26936 255320 26948
rect 255372 26936 255378 26988
rect 341058 26936 341064 26988
rect 341116 26976 341122 26988
rect 433334 26976 433340 26988
rect 341116 26948 433340 26976
rect 341116 26936 341122 26948
rect 433334 26936 433340 26948
rect 433392 26936 433398 26988
rect 77386 26868 77392 26920
rect 77444 26908 77450 26920
rect 218330 26908 218336 26920
rect 77444 26880 218336 26908
rect 77444 26868 77450 26880
rect 218330 26868 218336 26880
rect 218388 26868 218394 26920
rect 305178 26868 305184 26920
rect 305236 26908 305242 26920
rect 329834 26908 329840 26920
rect 305236 26880 329840 26908
rect 305236 26868 305242 26880
rect 329834 26868 329840 26880
rect 329892 26868 329898 26920
rect 385034 26868 385040 26920
rect 385092 26908 385098 26920
rect 564526 26908 564532 26920
rect 385092 26880 564532 26908
rect 385092 26868 385098 26880
rect 564526 26868 564532 26880
rect 564584 26868 564590 26920
rect 176746 25576 176752 25628
rect 176804 25616 176810 25628
rect 252830 25616 252836 25628
rect 176804 25588 252836 25616
rect 176804 25576 176810 25588
rect 252830 25576 252836 25588
rect 252888 25576 252894 25628
rect 311158 25576 311164 25628
rect 311216 25616 311222 25628
rect 339678 25616 339684 25628
rect 311216 25588 339684 25616
rect 311216 25576 311222 25588
rect 339678 25576 339684 25588
rect 339736 25576 339742 25628
rect 85666 25508 85672 25560
rect 85724 25548 85730 25560
rect 220906 25548 220912 25560
rect 85724 25520 220912 25548
rect 85724 25508 85730 25520
rect 220906 25508 220912 25520
rect 220964 25508 220970 25560
rect 258074 25508 258080 25560
rect 258132 25548 258138 25560
rect 280246 25548 280252 25560
rect 258132 25520 280252 25548
rect 258132 25508 258138 25520
rect 280246 25508 280252 25520
rect 280304 25508 280310 25560
rect 325694 25508 325700 25560
rect 325752 25548 325758 25560
rect 390830 25548 390836 25560
rect 325752 25520 390836 25548
rect 325752 25508 325758 25520
rect 390830 25508 390836 25520
rect 390888 25508 390894 25560
rect 392670 25508 392676 25560
rect 392728 25548 392734 25560
rect 568574 25548 568580 25560
rect 392728 25520 568580 25548
rect 392728 25508 392734 25520
rect 568574 25508 568580 25520
rect 568632 25508 568638 25560
rect 323026 24148 323032 24200
rect 323084 24188 323090 24200
rect 383654 24188 383660 24200
rect 323084 24160 383660 24188
rect 323084 24148 323090 24160
rect 383654 24148 383660 24160
rect 383712 24148 383718 24200
rect 172514 24080 172520 24132
rect 172572 24120 172578 24132
rect 251266 24120 251272 24132
rect 172572 24092 251272 24120
rect 172572 24080 172578 24092
rect 251266 24080 251272 24092
rect 251324 24080 251330 24132
rect 261110 24080 261116 24132
rect 261168 24120 261174 24132
rect 281810 24120 281816 24132
rect 261168 24092 281816 24120
rect 261168 24080 261174 24092
rect 281810 24080 281816 24092
rect 281868 24080 281874 24132
rect 382366 24080 382372 24132
rect 382424 24120 382430 24132
rect 554774 24120 554780 24132
rect 382424 24092 554780 24120
rect 382424 24080 382430 24092
rect 554774 24080 554780 24092
rect 554832 24080 554838 24132
rect 314654 22788 314660 22840
rect 314712 22828 314718 22840
rect 358814 22828 358820 22840
rect 314712 22800 358820 22828
rect 314712 22788 314718 22800
rect 358814 22788 358820 22800
rect 358872 22788 358878 22840
rect 168374 22720 168380 22772
rect 168432 22760 168438 22772
rect 249978 22760 249984 22772
rect 168432 22732 249984 22760
rect 168432 22720 168438 22732
rect 249978 22720 249984 22732
rect 250036 22720 250042 22772
rect 252554 22720 252560 22772
rect 252612 22760 252618 22772
rect 278958 22760 278964 22772
rect 252612 22732 278964 22760
rect 252612 22720 252618 22732
rect 278958 22720 278964 22732
rect 279016 22720 279022 22772
rect 298186 22720 298192 22772
rect 298244 22760 298250 22772
rect 310606 22760 310612 22772
rect 298244 22732 310612 22760
rect 298244 22720 298250 22732
rect 310606 22720 310612 22732
rect 310664 22720 310670 22772
rect 327074 22720 327080 22772
rect 327132 22760 327138 22772
rect 393314 22760 393320 22772
rect 327132 22732 393320 22760
rect 327132 22720 327138 22732
rect 393314 22720 393320 22732
rect 393372 22720 393378 22772
rect 396718 22720 396724 22772
rect 396776 22760 396782 22772
rect 550634 22760 550640 22772
rect 396776 22732 550640 22760
rect 396776 22720 396782 22732
rect 550634 22720 550640 22732
rect 550692 22720 550698 22772
rect 302326 21564 302332 21616
rect 302384 21604 302390 21616
rect 321646 21604 321652 21616
rect 302384 21576 321652 21604
rect 302384 21564 302390 21576
rect 321646 21564 321652 21576
rect 321704 21564 321710 21616
rect 321554 21428 321560 21480
rect 321612 21468 321618 21480
rect 378318 21468 378324 21480
rect 321612 21440 378324 21468
rect 321612 21428 321618 21440
rect 378318 21428 378324 21440
rect 378376 21428 378382 21480
rect 55214 21360 55220 21412
rect 55272 21400 55278 21412
rect 211430 21400 211436 21412
rect 55272 21372 211436 21400
rect 55272 21360 55278 21372
rect 211430 21360 211436 21372
rect 211488 21360 211494 21412
rect 214006 21360 214012 21412
rect 214064 21400 214070 21412
rect 265158 21400 265164 21412
rect 214064 21372 265164 21400
rect 214064 21360 214070 21372
rect 265158 21360 265164 21372
rect 265216 21360 265222 21412
rect 371326 21360 371332 21412
rect 371384 21400 371390 21412
rect 523126 21400 523132 21412
rect 371384 21372 523132 21400
rect 371384 21360 371390 21372
rect 523126 21360 523132 21372
rect 523184 21360 523190 21412
rect 393958 20612 393964 20664
rect 394016 20652 394022 20664
rect 580166 20652 580172 20664
rect 394016 20624 580172 20652
rect 394016 20612 394022 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 210050 20000 210056 20052
rect 210108 20040 210114 20052
rect 250438 20040 250444 20052
rect 210108 20012 250444 20040
rect 210108 20000 210114 20012
rect 250438 20000 250444 20012
rect 250496 20000 250502 20052
rect 319438 20000 319444 20052
rect 319496 20040 319502 20052
rect 363046 20040 363052 20052
rect 319496 20012 363052 20040
rect 319496 20000 319502 20012
rect 363046 20000 363052 20012
rect 363104 20000 363110 20052
rect 192110 19932 192116 19984
rect 192168 19972 192174 19984
rect 256878 19972 256884 19984
rect 192168 19944 256884 19972
rect 192168 19932 192174 19944
rect 256878 19932 256884 19944
rect 256936 19932 256942 19984
rect 334066 19932 334072 19984
rect 334124 19972 334130 19984
rect 415486 19972 415492 19984
rect 334124 19944 415492 19972
rect 334124 19932 334130 19944
rect 415486 19932 415492 19944
rect 415544 19932 415550 19984
rect 203058 18640 203064 18692
rect 203116 18680 203122 18692
rect 261018 18680 261024 18692
rect 203116 18652 261024 18680
rect 203116 18640 203122 18652
rect 261018 18640 261024 18652
rect 261076 18640 261082 18692
rect 309870 18640 309876 18692
rect 309928 18680 309934 18692
rect 338298 18680 338304 18692
rect 309928 18652 338304 18680
rect 309928 18640 309934 18652
rect 338298 18640 338304 18652
rect 338356 18640 338362 18692
rect 69106 18572 69112 18624
rect 69164 18612 69170 18624
rect 214558 18612 214564 18624
rect 69164 18584 214564 18612
rect 69164 18572 69170 18584
rect 214558 18572 214564 18584
rect 214616 18572 214622 18624
rect 263778 18572 263784 18624
rect 263836 18612 263842 18624
rect 281718 18612 281724 18624
rect 263836 18584 281724 18612
rect 263836 18572 263842 18584
rect 281718 18572 281724 18584
rect 281776 18572 281782 18624
rect 327810 18572 327816 18624
rect 327868 18612 327874 18624
rect 390922 18612 390928 18624
rect 327868 18584 390928 18612
rect 327868 18572 327874 18584
rect 390922 18572 390928 18584
rect 390980 18572 390986 18624
rect 392578 18572 392584 18624
rect 392636 18612 392642 18624
rect 518894 18612 518900 18624
rect 392636 18584 518900 18612
rect 392636 18572 392642 18584
rect 518894 18572 518900 18584
rect 518952 18572 518958 18624
rect 200390 17280 200396 17332
rect 200448 17320 200454 17332
rect 259546 17320 259552 17332
rect 200448 17292 259552 17320
rect 200448 17280 200454 17292
rect 259546 17280 259552 17292
rect 259604 17280 259610 17332
rect 315298 17280 315304 17332
rect 315356 17320 315362 17332
rect 323026 17320 323032 17332
rect 315356 17292 323032 17320
rect 315356 17280 315362 17292
rect 323026 17280 323032 17292
rect 323084 17280 323090 17332
rect 323578 17280 323584 17332
rect 323636 17320 323642 17332
rect 377030 17320 377036 17332
rect 323636 17292 377036 17320
rect 323636 17280 323642 17292
rect 377030 17280 377036 17292
rect 377088 17280 377094 17332
rect 37274 17212 37280 17264
rect 37332 17252 37338 17264
rect 203518 17252 203524 17264
rect 37332 17224 203524 17252
rect 37332 17212 37338 17224
rect 203518 17212 203524 17224
rect 203576 17212 203582 17264
rect 218054 17212 218060 17264
rect 218112 17252 218118 17264
rect 266630 17252 266636 17264
rect 218112 17224 266636 17252
rect 218112 17212 218118 17224
rect 266630 17212 266636 17224
rect 266688 17212 266694 17264
rect 301130 17212 301136 17264
rect 301188 17252 301194 17264
rect 317598 17252 317604 17264
rect 301188 17224 317604 17252
rect 301188 17212 301194 17224
rect 317598 17212 317604 17224
rect 317656 17212 317662 17264
rect 362954 17212 362960 17264
rect 363012 17252 363018 17264
rect 500954 17252 500960 17264
rect 363012 17224 500960 17252
rect 363012 17212 363018 17224
rect 500954 17212 500960 17224
rect 501012 17212 501018 17264
rect 211706 15920 211712 15972
rect 211764 15960 211770 15972
rect 263686 15960 263692 15972
rect 211764 15932 263692 15960
rect 211764 15920 211770 15932
rect 263686 15920 263692 15932
rect 263744 15920 263750 15972
rect 303798 15920 303804 15972
rect 303856 15960 303862 15972
rect 326338 15960 326344 15972
rect 303856 15932 326344 15960
rect 303856 15920 303862 15932
rect 326338 15920 326344 15932
rect 326396 15920 326402 15972
rect 51074 15852 51080 15904
rect 51132 15892 51138 15904
rect 188338 15892 188344 15904
rect 51132 15864 188344 15892
rect 51132 15852 51138 15864
rect 188338 15852 188344 15864
rect 188396 15852 188402 15904
rect 196802 15852 196808 15904
rect 196860 15892 196866 15904
rect 251818 15892 251824 15904
rect 196860 15864 251824 15892
rect 196860 15852 196866 15864
rect 251818 15852 251824 15864
rect 251876 15852 251882 15904
rect 256694 15852 256700 15904
rect 256752 15892 256758 15904
rect 273898 15892 273904 15904
rect 256752 15864 273904 15892
rect 256752 15852 256758 15864
rect 273898 15852 273904 15864
rect 273956 15852 273962 15904
rect 313366 15852 313372 15904
rect 313424 15892 313430 15904
rect 356330 15892 356336 15904
rect 313424 15864 356336 15892
rect 313424 15852 313430 15864
rect 356330 15852 356336 15864
rect 356388 15852 356394 15904
rect 368474 15852 368480 15904
rect 368532 15892 368538 15904
rect 515490 15892 515496 15904
rect 368532 15864 515496 15892
rect 368532 15852 368538 15864
rect 515490 15852 515496 15864
rect 515548 15852 515554 15904
rect 306466 14560 306472 14612
rect 306524 14600 306530 14612
rect 333882 14600 333888 14612
rect 306524 14572 333888 14600
rect 306524 14560 306530 14572
rect 333882 14560 333888 14572
rect 333940 14560 333946 14612
rect 221090 14492 221096 14544
rect 221148 14532 221154 14544
rect 267826 14532 267832 14544
rect 221148 14504 267832 14532
rect 221148 14492 221154 14504
rect 267826 14492 267832 14504
rect 267884 14492 267890 14544
rect 327718 14492 327724 14544
rect 327776 14532 327782 14544
rect 372890 14532 372896 14544
rect 327776 14504 372896 14532
rect 327776 14492 327782 14504
rect 372890 14492 372896 14504
rect 372948 14492 372954 14544
rect 168466 14424 168472 14476
rect 168524 14464 168530 14476
rect 235350 14464 235356 14476
rect 168524 14436 235356 14464
rect 168524 14424 168530 14436
rect 235350 14424 235356 14436
rect 235408 14424 235414 14476
rect 306558 14424 306564 14476
rect 306616 14464 306622 14476
rect 334618 14464 334624 14476
rect 306616 14436 334624 14464
rect 306616 14424 306622 14436
rect 334618 14424 334624 14436
rect 334676 14424 334682 14476
rect 364426 14424 364432 14476
rect 364484 14464 364490 14476
rect 505370 14464 505376 14476
rect 364484 14436 505376 14464
rect 364484 14424 364490 14436
rect 505370 14424 505376 14436
rect 505428 14424 505434 14476
rect 123018 13336 123024 13388
rect 123076 13376 123082 13388
rect 233326 13376 233332 13388
rect 123076 13348 233332 13376
rect 123076 13336 123082 13348
rect 233326 13336 233332 13348
rect 233384 13336 233390 13388
rect 119890 13268 119896 13320
rect 119948 13308 119954 13320
rect 231946 13308 231952 13320
rect 119948 13280 231952 13308
rect 119948 13268 119954 13280
rect 231946 13268 231952 13280
rect 232004 13268 232010 13320
rect 116394 13200 116400 13252
rect 116452 13240 116458 13252
rect 232130 13240 232136 13252
rect 116452 13212 232136 13240
rect 116452 13200 116458 13212
rect 232130 13200 232136 13212
rect 232188 13200 232194 13252
rect 367186 13200 367192 13252
rect 367244 13240 367250 13252
rect 511258 13240 511264 13252
rect 367244 13212 511264 13240
rect 367244 13200 367250 13212
rect 511258 13200 511264 13212
rect 511316 13200 511322 13252
rect 112346 13132 112352 13184
rect 112404 13172 112410 13184
rect 230566 13172 230572 13184
rect 112404 13144 230572 13172
rect 112404 13132 112410 13144
rect 230566 13132 230572 13144
rect 230624 13132 230630 13184
rect 303706 13132 303712 13184
rect 303764 13172 303770 13184
rect 327994 13172 328000 13184
rect 303764 13144 328000 13172
rect 303764 13132 303770 13144
rect 327994 13132 328000 13144
rect 328052 13132 328058 13184
rect 371234 13132 371240 13184
rect 371292 13172 371298 13184
rect 525426 13172 525432 13184
rect 371292 13144 525432 13172
rect 371292 13132 371298 13144
rect 525426 13132 525432 13144
rect 525484 13132 525490 13184
rect 22554 13064 22560 13116
rect 22612 13104 22618 13116
rect 198918 13104 198924 13116
rect 22612 13076 198924 13104
rect 22612 13064 22618 13076
rect 198918 13064 198924 13076
rect 198976 13064 198982 13116
rect 232038 13064 232044 13116
rect 232096 13104 232102 13116
rect 270678 13104 270684 13116
rect 232096 13076 270684 13104
rect 232096 13064 232102 13076
rect 270678 13064 270684 13076
rect 270736 13064 270742 13116
rect 270770 13064 270776 13116
rect 270828 13104 270834 13116
rect 284570 13104 284576 13116
rect 270828 13076 284576 13104
rect 270828 13064 270834 13076
rect 284570 13064 284576 13076
rect 284628 13064 284634 13116
rect 317506 13064 317512 13116
rect 317564 13104 317570 13116
rect 365714 13104 365720 13116
rect 317564 13076 365720 13104
rect 317564 13064 317570 13076
rect 365714 13064 365720 13076
rect 365772 13064 365778 13116
rect 374178 13064 374184 13116
rect 374236 13104 374242 13116
rect 532050 13104 532056 13116
rect 374236 13076 532056 13104
rect 374236 13064 374242 13076
rect 532050 13064 532056 13076
rect 532108 13064 532114 13116
rect 109034 12044 109040 12096
rect 109092 12084 109098 12096
rect 229186 12084 229192 12096
rect 109092 12056 229192 12084
rect 109092 12044 109098 12056
rect 229186 12044 229192 12056
rect 229244 12044 229250 12096
rect 105722 11976 105728 12028
rect 105780 12016 105786 12028
rect 227898 12016 227904 12028
rect 105780 11988 227904 12016
rect 105780 11976 105786 11988
rect 227898 11976 227904 11988
rect 227956 11976 227962 12028
rect 98178 11908 98184 11960
rect 98236 11948 98242 11960
rect 225046 11948 225052 11960
rect 98236 11920 225052 11948
rect 98236 11908 98242 11920
rect 225046 11908 225052 11920
rect 225104 11908 225110 11960
rect 93854 11840 93860 11892
rect 93912 11880 93918 11892
rect 223758 11880 223764 11892
rect 93912 11852 223764 11880
rect 93912 11840 93918 11852
rect 223758 11840 223764 11852
rect 223816 11840 223822 11892
rect 354858 11840 354864 11892
rect 354916 11880 354922 11892
rect 474090 11880 474096 11892
rect 354916 11852 474096 11880
rect 354916 11840 354922 11852
rect 474090 11840 474096 11852
rect 474148 11840 474154 11892
rect 84194 11772 84200 11824
rect 84252 11812 84258 11824
rect 220814 11812 220820 11824
rect 84252 11784 220820 11812
rect 84252 11772 84258 11784
rect 220814 11772 220820 11784
rect 220872 11772 220878 11824
rect 240134 11772 240140 11824
rect 240192 11812 240198 11824
rect 273346 11812 273352 11824
rect 240192 11784 273352 11812
rect 240192 11772 240198 11784
rect 273346 11772 273352 11784
rect 273404 11772 273410 11824
rect 301038 11772 301044 11824
rect 301096 11812 301102 11824
rect 320450 11812 320456 11824
rect 301096 11784 320456 11812
rect 301096 11772 301102 11784
rect 320450 11772 320456 11784
rect 320508 11772 320514 11824
rect 360378 11772 360384 11824
rect 360436 11812 360442 11824
rect 493042 11812 493048 11824
rect 360436 11784 493048 11812
rect 360436 11772 360442 11784
rect 493042 11772 493048 11784
rect 493100 11772 493106 11824
rect 80882 11704 80888 11756
rect 80940 11744 80946 11756
rect 219526 11744 219532 11756
rect 80940 11716 219532 11744
rect 80940 11704 80946 11716
rect 219526 11704 219532 11716
rect 219584 11704 219590 11756
rect 228266 11704 228272 11756
rect 228324 11744 228330 11756
rect 269758 11744 269764 11756
rect 228324 11716 269764 11744
rect 228324 11704 228330 11716
rect 269758 11704 269764 11716
rect 269816 11704 269822 11756
rect 310514 11704 310520 11756
rect 310572 11744 310578 11756
rect 349338 11744 349344 11756
rect 310572 11716 349344 11744
rect 310572 11704 310578 11716
rect 349338 11704 349344 11716
rect 349396 11704 349402 11756
rect 364334 11704 364340 11756
rect 364392 11744 364398 11756
rect 503714 11744 503720 11756
rect 364392 11716 503720 11744
rect 364392 11704 364398 11716
rect 503714 11704 503720 11716
rect 503772 11704 503778 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 168374 11636 168380 11688
rect 168432 11676 168438 11688
rect 169570 11676 169576 11688
rect 168432 11648 169576 11676
rect 168432 11636 168438 11648
rect 169570 11636 169576 11648
rect 169628 11636 169634 11688
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 331214 10820 331220 10872
rect 331272 10860 331278 10872
rect 407206 10860 407212 10872
rect 331272 10832 407212 10860
rect 331272 10820 331278 10832
rect 407206 10820 407212 10832
rect 407264 10820 407270 10872
rect 332686 10752 332692 10804
rect 332744 10792 332750 10804
rect 410794 10792 410800 10804
rect 332744 10764 410800 10792
rect 332744 10752 332750 10764
rect 410794 10752 410800 10764
rect 410852 10752 410858 10804
rect 333974 10684 333980 10736
rect 334032 10724 334038 10736
rect 414290 10724 414296 10736
rect 334032 10696 414296 10724
rect 334032 10684 334038 10696
rect 414290 10684 414296 10696
rect 414348 10684 414354 10736
rect 108114 10616 108120 10668
rect 108172 10656 108178 10668
rect 229370 10656 229376 10668
rect 108172 10628 229376 10656
rect 108172 10616 108178 10628
rect 229370 10616 229376 10628
rect 229428 10616 229434 10668
rect 335446 10616 335452 10668
rect 335504 10656 335510 10668
rect 417418 10656 417424 10668
rect 335504 10628 417424 10656
rect 335504 10616 335510 10628
rect 417418 10616 417424 10628
rect 417476 10616 417482 10668
rect 104066 10548 104072 10600
rect 104124 10588 104130 10600
rect 227806 10588 227812 10600
rect 104124 10560 227812 10588
rect 104124 10548 104130 10560
rect 227806 10548 227812 10560
rect 227864 10548 227870 10600
rect 335538 10548 335544 10600
rect 335596 10588 335602 10600
rect 420914 10588 420920 10600
rect 335596 10560 420920 10588
rect 335596 10548 335602 10560
rect 420914 10548 420920 10560
rect 420972 10548 420978 10600
rect 97442 10480 97448 10532
rect 97500 10520 97506 10532
rect 224954 10520 224960 10532
rect 97500 10492 224960 10520
rect 97500 10480 97506 10492
rect 224954 10480 224960 10492
rect 225012 10480 225018 10532
rect 336826 10480 336832 10532
rect 336884 10520 336890 10532
rect 423674 10520 423680 10532
rect 336884 10492 423680 10520
rect 336884 10480 336890 10492
rect 423674 10480 423680 10492
rect 423732 10480 423738 10532
rect 93946 10412 93952 10464
rect 94004 10452 94010 10464
rect 223666 10452 223672 10464
rect 94004 10424 223672 10452
rect 94004 10412 94010 10424
rect 223666 10412 223672 10424
rect 223724 10412 223730 10464
rect 267734 10412 267740 10464
rect 267792 10452 267798 10464
rect 283098 10452 283104 10464
rect 267792 10424 283104 10452
rect 267792 10412 267798 10424
rect 283098 10412 283104 10424
rect 283156 10412 283162 10464
rect 338206 10412 338212 10464
rect 338264 10452 338270 10464
rect 428458 10452 428464 10464
rect 338264 10424 428464 10452
rect 338264 10412 338270 10424
rect 428458 10412 428464 10424
rect 428516 10412 428522 10464
rect 52546 10344 52552 10396
rect 52604 10384 52610 10396
rect 209866 10384 209872 10396
rect 52604 10356 209872 10384
rect 52604 10344 52610 10356
rect 209866 10344 209872 10356
rect 209924 10344 209930 10396
rect 226334 10344 226340 10396
rect 226392 10384 226398 10396
rect 269206 10384 269212 10396
rect 226392 10356 269212 10384
rect 226392 10344 226398 10356
rect 269206 10344 269212 10356
rect 269264 10344 269270 10396
rect 302234 10344 302240 10396
rect 302292 10384 302298 10396
rect 324406 10384 324412 10396
rect 302292 10356 324412 10384
rect 302292 10344 302298 10356
rect 324406 10344 324412 10356
rect 324464 10344 324470 10396
rect 339586 10344 339592 10396
rect 339644 10384 339650 10396
rect 432046 10384 432052 10396
rect 339644 10356 432052 10384
rect 339644 10344 339650 10356
rect 432046 10344 432052 10356
rect 432104 10344 432110 10396
rect 44266 10276 44272 10328
rect 44324 10316 44330 10328
rect 207106 10316 207112 10328
rect 44324 10288 207112 10316
rect 44324 10276 44330 10288
rect 207106 10276 207112 10288
rect 207164 10276 207170 10328
rect 225138 10276 225144 10328
rect 225196 10316 225202 10328
rect 268378 10316 268384 10328
rect 225196 10288 268384 10316
rect 225196 10276 225202 10288
rect 268378 10276 268384 10288
rect 268436 10276 268442 10328
rect 305086 10276 305092 10328
rect 305144 10316 305150 10328
rect 332686 10316 332692 10328
rect 305144 10288 332692 10316
rect 305144 10276 305150 10288
rect 332686 10276 332692 10288
rect 332744 10276 332750 10328
rect 342346 10276 342352 10328
rect 342404 10316 342410 10328
rect 439130 10316 439136 10328
rect 342404 10288 439136 10316
rect 342404 10276 342410 10288
rect 439130 10276 439136 10288
rect 439188 10276 439194 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 309778 9596 309784 9648
rect 309836 9636 309842 9648
rect 315022 9636 315028 9648
rect 309836 9608 315028 9636
rect 309836 9596 309842 9608
rect 315022 9596 315028 9608
rect 315080 9596 315086 9648
rect 322934 9392 322940 9444
rect 322992 9432 322998 9444
rect 382366 9432 382372 9444
rect 322992 9404 382372 9432
rect 322992 9392 322998 9404
rect 382366 9392 382372 9404
rect 382424 9392 382430 9444
rect 372798 9324 372804 9376
rect 372856 9364 372862 9376
rect 527818 9364 527824 9376
rect 372856 9336 527824 9364
rect 372856 9324 372862 9336
rect 527818 9324 527824 9336
rect 527876 9324 527882 9376
rect 374086 9256 374092 9308
rect 374144 9296 374150 9308
rect 531314 9296 531320 9308
rect 374144 9268 531320 9296
rect 374144 9256 374150 9268
rect 531314 9256 531320 9268
rect 531372 9256 531378 9308
rect 376846 9188 376852 9240
rect 376904 9228 376910 9240
rect 538398 9228 538404 9240
rect 376904 9200 538404 9228
rect 376904 9188 376910 9200
rect 538398 9188 538404 9200
rect 538456 9188 538462 9240
rect 376938 9120 376944 9172
rect 376996 9160 377002 9172
rect 541986 9160 541992 9172
rect 376996 9132 541992 9160
rect 376996 9120 377002 9132
rect 541986 9120 541992 9132
rect 542044 9120 542050 9172
rect 239306 9052 239312 9104
rect 239364 9092 239370 9104
rect 265618 9092 265624 9104
rect 239364 9064 265624 9092
rect 239364 9052 239370 9064
rect 265618 9052 265624 9064
rect 265676 9052 265682 9104
rect 317414 9052 317420 9104
rect 317472 9092 317478 9104
rect 368198 9092 368204 9104
rect 317472 9064 368204 9092
rect 317472 9052 317478 9064
rect 368198 9052 368204 9064
rect 368256 9052 368262 9104
rect 378226 9052 378232 9104
rect 378284 9092 378290 9104
rect 545482 9092 545488 9104
rect 378284 9064 545488 9092
rect 378284 9052 378290 9064
rect 545482 9052 545488 9064
rect 545540 9052 545546 9104
rect 40678 8984 40684 9036
rect 40736 9024 40742 9036
rect 205726 9024 205732 9036
rect 40736 8996 205732 9024
rect 40736 8984 40742 8996
rect 205726 8984 205732 8996
rect 205784 8984 205790 9036
rect 208578 8984 208584 9036
rect 208636 9024 208642 9036
rect 263870 9024 263876 9036
rect 208636 8996 263876 9024
rect 208636 8984 208642 8996
rect 263870 8984 263876 8996
rect 263928 8984 263934 9036
rect 302878 8984 302884 9036
rect 302936 9024 302942 9036
rect 302936 8996 306374 9024
rect 302936 8984 302942 8996
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 196066 8956 196072 8968
rect 13596 8928 196072 8956
rect 13596 8916 13602 8928
rect 196066 8916 196072 8928
rect 196124 8916 196130 8968
rect 202690 8916 202696 8968
rect 202748 8956 202754 8968
rect 260926 8956 260932 8968
rect 202748 8928 260932 8956
rect 202748 8916 202754 8928
rect 260926 8916 260932 8928
rect 260984 8916 260990 8968
rect 295518 8916 295524 8968
rect 295576 8956 295582 8968
rect 303154 8956 303160 8968
rect 295576 8928 303160 8956
rect 295576 8916 295582 8928
rect 303154 8916 303160 8928
rect 303212 8916 303218 8968
rect 306346 8956 306374 8996
rect 318886 8984 318892 9036
rect 318944 9024 318950 9036
rect 371694 9024 371700 9036
rect 318944 8996 371700 9024
rect 318944 8984 318950 8996
rect 371694 8984 371700 8996
rect 371752 8984 371758 9036
rect 380894 8984 380900 9036
rect 380952 9024 380958 9036
rect 552658 9024 552664 9036
rect 380952 8996 552664 9024
rect 380952 8984 380958 8996
rect 552658 8984 552664 8996
rect 552716 8984 552722 9036
rect 310238 8956 310244 8968
rect 306346 8928 310244 8956
rect 310238 8916 310244 8928
rect 310296 8916 310302 8968
rect 320266 8916 320272 8968
rect 320324 8956 320330 8968
rect 375282 8956 375288 8968
rect 320324 8928 375288 8956
rect 320324 8916 320330 8928
rect 375282 8916 375288 8928
rect 375340 8916 375346 8968
rect 382274 8916 382280 8968
rect 382332 8956 382338 8968
rect 556154 8956 556160 8968
rect 382332 8928 556160 8956
rect 382332 8916 382338 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 83274 7828 83280 7880
rect 83332 7868 83338 7880
rect 219434 7868 219440 7880
rect 83332 7840 219440 7868
rect 83332 7828 83338 7840
rect 219434 7828 219440 7840
rect 219492 7828 219498 7880
rect 33594 7760 33600 7812
rect 33652 7800 33658 7812
rect 202966 7800 202972 7812
rect 33652 7772 202972 7800
rect 33652 7760 33658 7772
rect 202966 7760 202972 7772
rect 203024 7760 203030 7812
rect 350626 7760 350632 7812
rect 350684 7800 350690 7812
rect 462774 7800 462780 7812
rect 350684 7772 462780 7800
rect 350684 7760 350690 7772
rect 462774 7760 462780 7772
rect 462832 7760 462838 7812
rect 26510 7692 26516 7744
rect 26568 7732 26574 7744
rect 200298 7732 200304 7744
rect 26568 7704 200304 7732
rect 26568 7692 26574 7704
rect 200298 7692 200304 7704
rect 200356 7692 200362 7744
rect 229830 7692 229836 7744
rect 229888 7732 229894 7744
rect 270586 7732 270592 7744
rect 229888 7704 270592 7732
rect 229888 7692 229894 7704
rect 270586 7692 270592 7704
rect 270644 7692 270650 7744
rect 299566 7692 299572 7744
rect 299624 7732 299630 7744
rect 313826 7732 313832 7744
rect 299624 7704 313832 7732
rect 299624 7692 299630 7704
rect 313826 7692 313832 7704
rect 313884 7692 313890 7744
rect 353386 7692 353392 7744
rect 353444 7732 353450 7744
rect 473446 7732 473452 7744
rect 353444 7704 473452 7732
rect 353444 7692 353450 7704
rect 473446 7692 473452 7704
rect 473504 7692 473510 7744
rect 21818 7624 21824 7676
rect 21876 7664 21882 7676
rect 198826 7664 198832 7676
rect 21876 7636 198832 7664
rect 21876 7624 21882 7636
rect 198826 7624 198832 7636
rect 198884 7624 198890 7676
rect 222746 7624 222752 7676
rect 222804 7664 222810 7676
rect 267918 7664 267924 7676
rect 222804 7636 267924 7664
rect 222804 7624 222810 7636
rect 267918 7624 267924 7636
rect 267976 7624 267982 7676
rect 304994 7624 305000 7676
rect 305052 7664 305058 7676
rect 331582 7664 331588 7676
rect 305052 7636 331588 7664
rect 305052 7624 305058 7636
rect 331582 7624 331588 7636
rect 331640 7624 331646 7676
rect 333238 7624 333244 7676
rect 333296 7664 333302 7676
rect 345750 7664 345756 7676
rect 333296 7636 345756 7664
rect 333296 7624 333302 7636
rect 345750 7624 345756 7636
rect 345808 7624 345814 7676
rect 354766 7624 354772 7676
rect 354824 7664 354830 7676
rect 476942 7664 476948 7676
rect 354824 7636 476948 7664
rect 354824 7624 354830 7636
rect 476942 7624 476948 7636
rect 477000 7624 477006 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 193306 7596 193312 7608
rect 4120 7568 193312 7596
rect 4120 7556 4126 7568
rect 193306 7556 193312 7568
rect 193364 7556 193370 7608
rect 213362 7556 213368 7608
rect 213420 7596 213426 7608
rect 264238 7596 264244 7608
rect 213420 7568 264244 7596
rect 213420 7556 213426 7568
rect 264238 7556 264244 7568
rect 264296 7556 264302 7608
rect 313274 7556 313280 7608
rect 313332 7596 313338 7608
rect 354030 7596 354036 7608
rect 313332 7568 354036 7596
rect 313332 7556 313338 7568
rect 354030 7556 354036 7568
rect 354088 7556 354094 7608
rect 360194 7556 360200 7608
rect 360252 7596 360258 7608
rect 492306 7596 492312 7608
rect 360252 7568 492312 7596
rect 360252 7556 360258 7568
rect 492306 7556 492312 7568
rect 492364 7556 492370 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 189718 6848 189724 6860
rect 3476 6820 189724 6848
rect 3476 6808 3482 6820
rect 189718 6808 189724 6820
rect 189776 6808 189782 6860
rect 246390 6400 246396 6452
rect 246448 6440 246454 6452
rect 276106 6440 276112 6452
rect 246448 6412 276112 6440
rect 246448 6400 246454 6412
rect 276106 6400 276112 6412
rect 276164 6400 276170 6452
rect 242986 6332 242992 6384
rect 243044 6372 243050 6384
rect 274910 6372 274916 6384
rect 243044 6344 274916 6372
rect 243044 6332 243050 6344
rect 274910 6332 274916 6344
rect 274968 6332 274974 6384
rect 309134 6332 309140 6384
rect 309192 6372 309198 6384
rect 343358 6372 343364 6384
rect 309192 6344 343364 6372
rect 309192 6332 309198 6344
rect 343358 6332 343364 6344
rect 343416 6332 343422 6384
rect 207382 6264 207388 6316
rect 207440 6304 207446 6316
rect 247678 6304 247684 6316
rect 207440 6276 247684 6304
rect 207440 6264 207446 6276
rect 247678 6264 247684 6276
rect 247736 6264 247742 6316
rect 332594 6264 332600 6316
rect 332652 6304 332658 6316
rect 413094 6304 413100 6316
rect 332652 6276 413100 6304
rect 332652 6264 332658 6276
rect 413094 6264 413100 6276
rect 413152 6264 413158 6316
rect 205082 6196 205088 6248
rect 205140 6236 205146 6248
rect 253198 6236 253204 6248
rect 205140 6208 253204 6236
rect 205140 6196 205146 6208
rect 253198 6196 253204 6208
rect 253256 6196 253262 6248
rect 300946 6196 300952 6248
rect 301004 6236 301010 6248
rect 317322 6236 317328 6248
rect 301004 6208 317328 6236
rect 301004 6196 301010 6208
rect 317322 6196 317328 6208
rect 317380 6196 317386 6248
rect 335354 6196 335360 6248
rect 335412 6236 335418 6248
rect 420178 6236 420184 6248
rect 335412 6208 420184 6236
rect 335412 6196 335418 6208
rect 420178 6196 420184 6208
rect 420236 6196 420242 6248
rect 65518 6128 65524 6180
rect 65576 6168 65582 6180
rect 214098 6168 214104 6180
rect 65576 6140 214104 6168
rect 65576 6128 65582 6140
rect 214098 6128 214104 6140
rect 214156 6128 214162 6180
rect 227530 6128 227536 6180
rect 227588 6168 227594 6180
rect 269298 6168 269304 6180
rect 227588 6140 269304 6168
rect 227588 6128 227594 6140
rect 269298 6128 269304 6140
rect 269356 6128 269362 6180
rect 303614 6128 303620 6180
rect 303672 6168 303678 6180
rect 325602 6168 325608 6180
rect 303672 6140 325608 6168
rect 303672 6128 303678 6140
rect 325602 6128 325608 6140
rect 325660 6128 325666 6180
rect 336734 6128 336740 6180
rect 336792 6168 336798 6180
rect 423766 6168 423772 6180
rect 336792 6140 423772 6168
rect 336792 6128 336798 6140
rect 423766 6128 423772 6140
rect 423824 6128 423830 6180
rect 390554 5176 390560 5228
rect 390612 5216 390618 5228
rect 390922 5216 390928 5228
rect 390612 5188 390928 5216
rect 390612 5176 390618 5188
rect 390922 5176 390928 5188
rect 390980 5176 390986 5228
rect 367094 5108 367100 5160
rect 367152 5148 367158 5160
rect 512454 5148 512460 5160
rect 367152 5120 512460 5148
rect 367152 5108 367158 5120
rect 512454 5108 512460 5120
rect 512512 5108 512518 5160
rect 54938 5040 54944 5092
rect 54996 5080 55002 5092
rect 209866 5080 209872 5092
rect 54996 5052 209872 5080
rect 54996 5040 55002 5052
rect 209866 5040 209872 5052
rect 209924 5040 209930 5092
rect 372706 5040 372712 5092
rect 372764 5080 372770 5092
rect 526622 5080 526628 5092
rect 372764 5052 526628 5080
rect 372764 5040 372770 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 195974 5012 195980 5024
rect 12400 4984 195980 5012
rect 12400 4972 12406 4984
rect 195974 4972 195980 4984
rect 196032 4972 196038 5024
rect 218146 4972 218152 5024
rect 218204 5012 218210 5024
rect 235258 5012 235264 5024
rect 218204 4984 235264 5012
rect 218204 4972 218210 4984
rect 235258 4972 235264 4984
rect 235316 4972 235322 5024
rect 249978 4972 249984 5024
rect 250036 5012 250042 5024
rect 277670 5012 277676 5024
rect 250036 4984 277676 5012
rect 250036 4972 250042 4984
rect 277670 4972 277676 4984
rect 277728 4972 277734 5024
rect 372614 4972 372620 5024
rect 372672 5012 372678 5024
rect 530118 5012 530124 5024
rect 372672 4984 530124 5012
rect 372672 4972 372678 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 191834 4944 191840 4956
rect 2924 4916 191840 4944
rect 2924 4904 2930 4916
rect 191834 4904 191840 4916
rect 191892 4904 191898 4956
rect 235810 4904 235816 4956
rect 235868 4944 235874 4956
rect 271966 4944 271972 4956
rect 235868 4916 271972 4944
rect 235868 4904 235874 4916
rect 271966 4904 271972 4916
rect 272024 4904 272030 4956
rect 306374 4904 306380 4956
rect 306432 4944 306438 4956
rect 336274 4944 336280 4956
rect 306432 4916 336280 4944
rect 306432 4904 306438 4916
rect 336274 4904 336280 4916
rect 336332 4904 336338 4956
rect 373994 4904 374000 4956
rect 374052 4944 374058 4956
rect 533706 4944 533712 4956
rect 374052 4916 533712 4944
rect 374052 4904 374058 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 192018 4876 192024 4888
rect 1728 4848 192024 4876
rect 1728 4836 1734 4848
rect 192018 4836 192024 4848
rect 192076 4836 192082 4888
rect 201494 4836 201500 4888
rect 201552 4876 201558 4888
rect 260834 4876 260840 4888
rect 201552 4848 260840 4876
rect 201552 4836 201558 4848
rect 260834 4836 260840 4848
rect 260892 4836 260898 4888
rect 318794 4836 318800 4888
rect 318852 4876 318858 4888
rect 370590 4876 370596 4888
rect 318852 4848 370596 4876
rect 318852 4836 318858 4848
rect 370590 4836 370596 4848
rect 370648 4836 370654 4888
rect 376754 4836 376760 4888
rect 376812 4876 376818 4888
rect 540790 4876 540796 4888
rect 376812 4848 540796 4876
rect 376812 4836 376818 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 191926 4808 191932 4820
rect 624 4780 191932 4808
rect 624 4768 630 4780
rect 191926 4768 191932 4780
rect 191984 4768 191990 4820
rect 195606 4768 195612 4820
rect 195664 4808 195670 4820
rect 257338 4808 257344 4820
rect 195664 4780 257344 4808
rect 195664 4768 195670 4780
rect 257338 4768 257344 4780
rect 257396 4768 257402 4820
rect 320174 4768 320180 4820
rect 320232 4808 320238 4820
rect 374086 4808 374092 4820
rect 320232 4780 374092 4808
rect 320232 4768 320238 4780
rect 374086 4768 374092 4780
rect 374144 4768 374150 4820
rect 378134 4768 378140 4820
rect 378192 4808 378198 4820
rect 544378 4808 544384 4820
rect 378192 4780 544384 4808
rect 378192 4768 378198 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 300118 4496 300124 4548
rect 300176 4536 300182 4548
rect 306742 4536 306748 4548
rect 300176 4508 306748 4536
rect 300176 4496 300182 4508
rect 306742 4496 306748 4508
rect 306800 4496 306806 4548
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 347038 4156 347044 4208
rect 347096 4196 347102 4208
rect 352834 4196 352840 4208
rect 347096 4168 352840 4196
rect 347096 4156 347102 4168
rect 352834 4156 352840 4168
rect 352892 4156 352898 4208
rect 46658 4088 46664 4140
rect 46716 4128 46722 4140
rect 207014 4128 207020 4140
rect 46716 4100 207020 4128
rect 46716 4088 46722 4100
rect 207014 4088 207020 4100
rect 207072 4088 207078 4140
rect 265342 4088 265348 4140
rect 265400 4128 265406 4140
rect 282914 4128 282920 4140
rect 265400 4100 282920 4128
rect 265400 4088 265406 4100
rect 282914 4088 282920 4100
rect 282972 4088 282978 4140
rect 285398 4088 285404 4140
rect 285456 4128 285462 4140
rect 289078 4128 289084 4140
rect 285456 4100 289084 4128
rect 285456 4088 285462 4100
rect 289078 4088 289084 4100
rect 289136 4088 289142 4140
rect 345014 4088 345020 4140
rect 345072 4128 345078 4140
rect 447410 4128 447416 4140
rect 345072 4100 447416 4128
rect 345072 4088 345078 4100
rect 447410 4088 447416 4100
rect 447468 4088 447474 4140
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 205634 4060 205640 4072
rect 43128 4032 205640 4060
rect 43128 4020 43134 4032
rect 205634 4020 205640 4032
rect 205692 4020 205698 4072
rect 262950 4020 262956 4072
rect 263008 4060 263014 4072
rect 281626 4060 281632 4072
rect 263008 4032 281632 4060
rect 263008 4020 263014 4032
rect 281626 4020 281632 4032
rect 281684 4020 281690 4072
rect 283098 4020 283104 4072
rect 283156 4060 283162 4072
rect 288526 4060 288532 4072
rect 283156 4032 288532 4060
rect 283156 4020 283162 4032
rect 288526 4020 288532 4032
rect 288584 4020 288590 4072
rect 347774 4020 347780 4072
rect 347832 4060 347838 4072
rect 454494 4060 454500 4072
rect 347832 4032 454500 4060
rect 347832 4020 347838 4032
rect 454494 4020 454500 4032
rect 454552 4020 454558 4072
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 204530 3992 204536 4004
rect 39632 3964 204536 3992
rect 39632 3952 39638 3964
rect 204530 3952 204536 3964
rect 204588 3952 204594 4004
rect 259546 3952 259552 4004
rect 259604 3992 259610 4004
rect 280338 3992 280344 4004
rect 259604 3964 280344 3992
rect 259604 3952 259610 3964
rect 280338 3952 280344 3964
rect 280396 3952 280402 4004
rect 280706 3952 280712 4004
rect 280764 3992 280770 4004
rect 287238 3992 287244 4004
rect 280764 3964 287244 3992
rect 280764 3952 280770 3964
rect 287238 3952 287244 3964
rect 287296 3952 287302 4004
rect 295978 3952 295984 4004
rect 296036 3992 296042 4004
rect 299658 3992 299664 4004
rect 296036 3964 299664 3992
rect 296036 3952 296042 3964
rect 299658 3952 299664 3964
rect 299716 3952 299722 4004
rect 349246 3952 349252 4004
rect 349304 3992 349310 4004
rect 458082 3992 458088 4004
rect 349304 3964 458088 3992
rect 349304 3952 349310 3964
rect 458082 3952 458088 3964
rect 458140 3952 458146 4004
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 204346 3924 204352 3936
rect 36044 3896 204352 3924
rect 36044 3884 36050 3896
rect 204346 3884 204352 3896
rect 204404 3884 204410 3936
rect 255866 3884 255872 3936
rect 255924 3924 255930 3936
rect 278866 3924 278872 3936
rect 255924 3896 278872 3924
rect 255924 3884 255930 3896
rect 278866 3884 278872 3896
rect 278924 3884 278930 3936
rect 295334 3884 295340 3936
rect 295392 3924 295398 3936
rect 301958 3924 301964 3936
rect 295392 3896 301964 3924
rect 295392 3884 295398 3896
rect 301958 3884 301964 3896
rect 302016 3884 302022 3936
rect 349154 3884 349160 3936
rect 349212 3924 349218 3936
rect 461578 3924 461584 3936
rect 349212 3896 461584 3924
rect 349212 3884 349218 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 32398 3816 32404 3868
rect 32456 3856 32462 3868
rect 202874 3856 202880 3868
rect 32456 3828 202880 3856
rect 32456 3816 32462 3828
rect 202874 3816 202880 3828
rect 202932 3816 202938 3868
rect 252370 3816 252376 3868
rect 252428 3856 252434 3868
rect 277578 3856 277584 3868
rect 252428 3828 277584 3856
rect 252428 3816 252434 3828
rect 277578 3816 277584 3828
rect 277636 3816 277642 3868
rect 350534 3816 350540 3868
rect 350592 3856 350598 3868
rect 465166 3856 465172 3868
rect 350592 3828 465172 3856
rect 350592 3816 350598 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 201770 3788 201776 3800
rect 28960 3760 201776 3788
rect 28960 3748 28966 3760
rect 201770 3748 201776 3760
rect 201828 3748 201834 3800
rect 248782 3748 248788 3800
rect 248840 3788 248846 3800
rect 277486 3788 277492 3800
rect 248840 3760 277492 3788
rect 248840 3748 248846 3760
rect 277486 3748 277492 3760
rect 277544 3748 277550 3800
rect 296806 3748 296812 3800
rect 296864 3788 296870 3800
rect 309042 3788 309048 3800
rect 296864 3760 309048 3788
rect 296864 3748 296870 3760
rect 309042 3748 309048 3760
rect 309100 3748 309106 3800
rect 351914 3748 351920 3800
rect 351972 3788 351978 3800
rect 468662 3788 468668 3800
rect 351972 3760 468668 3788
rect 351972 3748 351978 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 200206 3720 200212 3732
rect 25372 3692 200212 3720
rect 25372 3680 25378 3692
rect 200206 3680 200212 3692
rect 200264 3680 200270 3732
rect 245194 3680 245200 3732
rect 245252 3720 245258 3732
rect 276198 3720 276204 3732
rect 245252 3692 276204 3720
rect 245252 3680 245258 3692
rect 276198 3680 276204 3692
rect 276256 3680 276262 3732
rect 293954 3680 293960 3732
rect 294012 3720 294018 3732
rect 297266 3720 297272 3732
rect 294012 3692 297272 3720
rect 294012 3680 294018 3692
rect 297266 3680 297272 3692
rect 297324 3680 297330 3732
rect 297376 3692 306374 3720
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 21358 3652 21364 3664
rect 14792 3624 21364 3652
rect 14792 3612 14798 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 200114 3652 200120 3664
rect 24268 3624 200120 3652
rect 24268 3612 24274 3624
rect 200114 3612 200120 3624
rect 200172 3612 200178 3664
rect 241698 3612 241704 3664
rect 241756 3652 241762 3664
rect 274726 3652 274732 3664
rect 241756 3624 274732 3652
rect 241756 3612 241762 3624
rect 274726 3612 274732 3624
rect 274784 3612 274790 3664
rect 276014 3612 276020 3664
rect 276072 3652 276078 3664
rect 285858 3652 285864 3664
rect 276072 3624 285864 3652
rect 276072 3612 276078 3624
rect 285858 3612 285864 3624
rect 285916 3612 285922 3664
rect 296714 3612 296720 3664
rect 296772 3652 296778 3664
rect 297376 3652 297404 3692
rect 296772 3624 297404 3652
rect 296772 3612 296778 3624
rect 298094 3612 298100 3664
rect 298152 3652 298158 3664
rect 306346 3652 306374 3692
rect 353294 3680 353300 3732
rect 353352 3720 353358 3732
rect 472250 3720 472256 3732
rect 353352 3692 472256 3720
rect 353352 3680 353358 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 307938 3652 307944 3664
rect 298152 3624 304488 3652
rect 306346 3624 307944 3652
rect 298152 3612 298158 3624
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 197630 3584 197636 3596
rect 19484 3556 197636 3584
rect 19484 3544 19490 3556
rect 197630 3544 197636 3556
rect 197688 3544 197694 3596
rect 238110 3544 238116 3596
rect 238168 3584 238174 3596
rect 273530 3584 273536 3596
rect 238168 3556 273536 3584
rect 238168 3544 238174 3556
rect 273530 3544 273536 3556
rect 273588 3544 273594 3596
rect 277118 3544 277124 3596
rect 277176 3584 277182 3596
rect 287146 3584 287152 3596
rect 277176 3556 287152 3584
rect 277176 3544 277182 3556
rect 287146 3544 287152 3556
rect 287204 3544 287210 3596
rect 290182 3544 290188 3596
rect 290240 3584 290246 3596
rect 291286 3584 291292 3596
rect 290240 3556 291292 3584
rect 290240 3544 290246 3556
rect 291286 3544 291292 3556
rect 291344 3544 291350 3596
rect 292574 3544 292580 3596
rect 292632 3584 292638 3596
rect 293310 3584 293316 3596
rect 292632 3556 293316 3584
rect 292632 3544 292638 3556
rect 293310 3544 293316 3556
rect 293368 3544 293374 3596
rect 295426 3544 295432 3596
rect 295484 3584 295490 3596
rect 304350 3584 304356 3596
rect 295484 3556 304356 3584
rect 295484 3544 295490 3556
rect 304350 3544 304356 3556
rect 304408 3544 304414 3596
rect 304460 3584 304488 3624
rect 307938 3612 307944 3624
rect 307996 3612 308002 3664
rect 354674 3612 354680 3664
rect 354732 3652 354738 3664
rect 475746 3652 475752 3664
rect 354732 3624 475752 3652
rect 354732 3612 354738 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 312630 3584 312636 3596
rect 304460 3556 312636 3584
rect 312630 3544 312636 3556
rect 312688 3544 312694 3596
rect 356054 3544 356060 3596
rect 356112 3584 356118 3596
rect 356112 3556 364334 3584
rect 356112 3544 356118 3556
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 18598 3516 18604 3528
rect 17092 3488 18604 3516
rect 17092 3476 17098 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 198734 3516 198740 3528
rect 20680 3488 198740 3516
rect 20680 3476 20686 3488
rect 198734 3476 198740 3488
rect 198792 3476 198798 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219250 3516 219256 3528
rect 218112 3488 219256 3516
rect 218112 3476 218118 3488
rect 219250 3476 219256 3488
rect 219308 3476 219314 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260650 3516 260656 3528
rect 259512 3488 260656 3516
rect 259512 3476 259518 3488
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 272426 3476 272432 3528
rect 272484 3516 272490 3528
rect 284386 3516 284392 3528
rect 272484 3488 284392 3516
rect 272484 3476 272490 3488
rect 284386 3476 284392 3488
rect 284444 3476 284450 3528
rect 294046 3476 294052 3528
rect 294104 3516 294110 3528
rect 298462 3516 298468 3528
rect 294104 3488 298468 3516
rect 294104 3476 294110 3488
rect 298462 3476 298468 3488
rect 298520 3476 298526 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 316218 3516 316224 3528
rect 299532 3488 316224 3516
rect 299532 3476 299538 3488
rect 316218 3476 316224 3488
rect 316276 3476 316282 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 357526 3476 357532 3528
rect 357584 3516 357590 3528
rect 358722 3516 358728 3528
rect 357584 3488 358728 3516
rect 357584 3476 357590 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 364306 3516 364334 3556
rect 390738 3544 390744 3596
rect 390796 3584 390802 3596
rect 582190 3584 582196 3596
rect 390796 3556 582196 3584
rect 390796 3544 390802 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 479334 3516 479340 3528
rect 364306 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 547874 3476 547880 3528
rect 547932 3516 547938 3528
rect 548702 3516 548708 3528
rect 547932 3488 548708 3516
rect 547932 3476 547938 3488
rect 548702 3476 548708 3488
rect 548760 3476 548766 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 570598 3476 570604 3528
rect 570656 3516 570662 3528
rect 571518 3516 571524 3528
rect 570656 3488 571524 3516
rect 570656 3476 570662 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 572714 3516 572720 3528
rect 572036 3488 572720 3516
rect 572036 3476 572042 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 10318 3448 10324 3460
rect 6512 3420 10324 3448
rect 6512 3408 6518 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 17218 3448 17224 3460
rect 15988 3420 17224 3448
rect 15988 3408 15994 3420
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 194778 3448 194784 3460
rect 26206 3420 194784 3448
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 26206 3380 26234 3420
rect 194778 3408 194784 3420
rect 194836 3408 194842 3460
rect 231026 3408 231032 3460
rect 231084 3448 231090 3460
rect 270862 3448 270868 3460
rect 231084 3420 270868 3448
rect 231084 3408 231090 3420
rect 270862 3408 270868 3420
rect 270920 3408 270926 3460
rect 273622 3408 273628 3460
rect 273680 3448 273686 3460
rect 285766 3448 285772 3460
rect 273680 3420 285772 3448
rect 273680 3408 273686 3420
rect 285766 3408 285772 3420
rect 285824 3408 285830 3460
rect 300854 3408 300860 3460
rect 300912 3448 300918 3460
rect 319714 3448 319720 3460
rect 300912 3420 319720 3448
rect 300912 3408 300918 3420
rect 319714 3408 319720 3420
rect 319772 3408 319778 3460
rect 365714 3408 365720 3460
rect 365772 3448 365778 3460
rect 367002 3448 367008 3460
rect 365772 3420 367008 3448
rect 365772 3408 365778 3420
rect 367002 3408 367008 3420
rect 367060 3408 367066 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 580994 3448 581000 3460
rect 390612 3420 581000 3448
rect 390612 3408 390618 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 11204 3352 26234 3380
rect 11204 3340 11210 3352
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 227714 3380 227720 3392
rect 106976 3352 227720 3380
rect 106976 3340 106982 3352
rect 227714 3340 227720 3352
rect 227772 3340 227778 3392
rect 266538 3340 266544 3392
rect 266596 3380 266602 3392
rect 283006 3380 283012 3392
rect 266596 3352 283012 3380
rect 266596 3340 266602 3352
rect 283006 3340 283012 3352
rect 283064 3340 283070 3392
rect 296898 3340 296904 3392
rect 296956 3380 296962 3392
rect 305546 3380 305552 3392
rect 296956 3352 305552 3380
rect 296956 3340 296962 3352
rect 305546 3340 305552 3352
rect 305604 3340 305610 3392
rect 342254 3340 342260 3392
rect 342312 3380 342318 3392
rect 440234 3380 440240 3392
rect 342312 3352 440240 3380
rect 342312 3340 342318 3352
rect 440234 3340 440240 3352
rect 440292 3340 440298 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 572070 3340 572076 3392
rect 572128 3380 572134 3392
rect 573910 3380 573916 3392
rect 572128 3352 573916 3380
rect 572128 3340 572134 3352
rect 573910 3340 573916 3352
rect 573968 3340 573974 3392
rect 114002 3272 114008 3324
rect 114060 3312 114066 3324
rect 230474 3312 230480 3324
rect 114060 3284 230480 3312
rect 114060 3272 114066 3284
rect 230474 3272 230480 3284
rect 230532 3272 230538 3324
rect 268838 3272 268844 3324
rect 268896 3312 268902 3324
rect 284294 3312 284300 3324
rect 268896 3284 284300 3312
rect 268896 3272 268902 3284
rect 284294 3272 284300 3284
rect 284352 3272 284358 3324
rect 339494 3272 339500 3324
rect 339552 3312 339558 3324
rect 433242 3312 433248 3324
rect 339552 3284 433248 3312
rect 339552 3272 339558 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 121086 3204 121092 3256
rect 121144 3244 121150 3256
rect 233234 3244 233240 3256
rect 121144 3216 233240 3244
rect 121144 3204 121150 3216
rect 233234 3204 233240 3216
rect 233292 3204 233298 3256
rect 270034 3204 270040 3256
rect 270092 3244 270098 3256
rect 284478 3244 284484 3256
rect 270092 3216 284484 3244
rect 270092 3204 270098 3216
rect 284478 3204 284484 3216
rect 284536 3204 284542 3256
rect 297358 3204 297364 3256
rect 297416 3244 297422 3256
rect 300762 3244 300768 3256
rect 297416 3216 300768 3244
rect 297416 3204 297422 3216
rect 300762 3204 300768 3216
rect 300820 3204 300826 3256
rect 338114 3204 338120 3256
rect 338172 3244 338178 3256
rect 338172 3216 412634 3244
rect 338172 3204 338178 3216
rect 234614 3136 234620 3188
rect 234672 3176 234678 3188
rect 272058 3176 272064 3188
rect 234672 3148 272064 3176
rect 234672 3136 234678 3148
rect 272058 3136 272064 3148
rect 272116 3136 272122 3188
rect 292850 3136 292856 3188
rect 292908 3176 292914 3188
rect 296070 3176 296076 3188
rect 292908 3148 296076 3176
rect 292908 3136 292914 3148
rect 296070 3136 296076 3148
rect 296128 3136 296134 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 407114 3136 407120 3188
rect 407172 3176 407178 3188
rect 408402 3176 408408 3188
rect 407172 3148 408408 3176
rect 407172 3136 407178 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 412606 3176 412634 3216
rect 415394 3204 415400 3256
rect 415452 3244 415458 3256
rect 416682 3244 416688 3256
rect 415452 3216 416688 3244
rect 415452 3204 415458 3216
rect 416682 3204 416688 3216
rect 416740 3204 416746 3256
rect 423674 3204 423680 3256
rect 423732 3244 423738 3256
rect 424962 3244 424968 3256
rect 423732 3216 424968 3244
rect 423732 3204 423738 3216
rect 424962 3204 424968 3216
rect 425020 3204 425026 3256
rect 426158 3176 426164 3188
rect 412606 3148 426164 3176
rect 426158 3136 426164 3148
rect 426216 3136 426222 3188
rect 284294 3000 284300 3052
rect 284352 3040 284358 3052
rect 288618 3040 288624 3052
rect 284352 3012 288624 3040
rect 284352 3000 284358 3012
rect 288618 3000 288624 3012
rect 288676 3000 288682 3052
rect 292758 3000 292764 3052
rect 292816 3040 292822 3052
rect 294874 3040 294880 3052
rect 292816 3012 294880 3040
rect 292816 3000 292822 3012
rect 294874 3000 294880 3012
rect 294932 3000 294938 3052
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 14458 2904 14464 2916
rect 10008 2876 14464 2904
rect 10008 2864 10014 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 328460 700816 328512 700868
rect 397460 700816 397512 700868
rect 335360 700748 335412 700800
rect 413652 700748 413704 700800
rect 343640 700680 343692 700732
rect 429844 700680 429896 700732
rect 350540 700612 350592 700664
rect 462320 700612 462372 700664
rect 357440 700544 357492 700596
rect 478512 700544 478564 700596
rect 365720 700476 365772 700528
rect 494796 700476 494848 700528
rect 306380 700408 306432 700460
rect 332508 700408 332560 700460
rect 372620 700408 372672 700460
rect 527180 700408 527232 700460
rect 313280 700340 313332 700392
rect 348792 700340 348844 700392
rect 379520 700340 379572 700392
rect 543464 700340 543516 700392
rect 321560 700272 321612 700324
rect 364984 700272 365036 700324
rect 387800 700272 387852 700324
rect 559656 700272 559708 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 3424 683136 3476 683188
rect 18604 683136 18656 683188
rect 406384 683136 406436 683188
rect 579620 683136 579672 683188
rect 395344 670692 395396 670744
rect 580172 670692 580224 670744
rect 400864 643084 400916 643136
rect 580172 643084 580224 643136
rect 3332 632068 3384 632120
rect 21364 632068 21416 632120
rect 393964 630640 394016 630692
rect 579988 630640 580040 630692
rect 3332 618264 3384 618316
rect 13084 618264 13136 618316
rect 2780 605888 2832 605940
rect 4804 605888 4856 605940
rect 3332 579640 3384 579692
rect 22744 579640 22796 579692
rect 405004 576852 405056 576904
rect 579988 576852 580040 576904
rect 399484 536800 399536 536852
rect 579620 536800 579672 536852
rect 2964 527144 3016 527196
rect 26884 527144 26936 527196
rect 3332 514768 3384 514820
rect 14464 514768 14516 514820
rect 3332 501304 3384 501356
rect 8944 501304 8996 501356
rect 3332 474716 3384 474768
rect 32404 474716 32456 474768
rect 403624 470568 403676 470620
rect 579988 470568 580040 470620
rect 549904 456764 549956 456816
rect 580172 456764 580224 456816
rect 407764 418140 407816 418192
rect 580172 418140 580224 418192
rect 3332 409844 3384 409896
rect 17224 409844 17276 409896
rect 396724 404336 396776 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 10324 397468 10376 397520
rect 169760 393116 169812 393168
rect 254952 393116 255004 393168
rect 153200 393048 153252 393100
rect 247500 393048 247552 393100
rect 136640 392980 136692 393032
rect 240140 392980 240192 393032
rect 104900 392912 104952 392964
rect 232688 392912 232740 392964
rect 88340 392844 88392 392896
rect 225328 392844 225380 392896
rect 71780 392776 71832 392828
rect 217876 392776 217928 392828
rect 40040 392708 40092 392760
rect 210516 392708 210568 392760
rect 234620 392708 234672 392760
rect 277124 392708 277176 392760
rect 23480 392640 23532 392692
rect 203064 392640 203116 392692
rect 218060 392640 218112 392692
rect 269764 392640 269816 392692
rect 282920 392640 282972 392692
rect 291936 392640 291988 392692
rect 6920 392572 6972 392624
rect 195704 392572 195756 392624
rect 201500 392572 201552 392624
rect 262312 392572 262364 392624
rect 266360 392572 266412 392624
rect 284576 392572 284628 392624
rect 18604 387744 18656 387796
rect 189080 387744 189132 387796
rect 394516 387744 394568 387796
rect 580264 387744 580316 387796
rect 3424 380808 3476 380860
rect 189080 380808 189132 380860
rect 394608 380808 394660 380860
rect 406384 380808 406436 380860
rect 394148 375300 394200 375352
rect 395344 375300 395396 375352
rect 3516 373940 3568 373992
rect 189080 373940 189132 373992
rect 393872 368092 393924 368144
rect 400864 368092 400916 368144
rect 21364 367004 21416 367056
rect 189080 367004 189132 367056
rect 394056 364352 394108 364404
rect 580172 364352 580224 364404
rect 13084 360136 13136 360188
rect 189080 360136 189132 360188
rect 394608 355988 394660 356040
rect 580356 355988 580408 356040
rect 4804 353200 4856 353252
rect 189080 353200 189132 353252
rect 394608 350480 394660 350532
rect 580448 350480 580500 350532
rect 22744 347692 22796 347744
rect 189080 347692 189132 347744
rect 394240 343544 394292 343596
rect 405004 343544 405056 343596
rect 3608 340824 3660 340876
rect 189080 340824 189132 340876
rect 394608 338036 394660 338088
rect 580540 338036 580592 338088
rect 3700 333888 3752 333940
rect 189080 333888 189132 333940
rect 393964 331168 394016 331220
rect 399484 331168 399536 331220
rect 26884 327020 26936 327072
rect 189080 327020 189132 327072
rect 394608 325592 394660 325644
rect 580632 325592 580684 325644
rect 14464 320084 14516 320136
rect 189080 320084 189132 320136
rect 394608 318724 394660 318776
rect 580724 318724 580776 318776
rect 8944 314576 8996 314628
rect 189080 314576 189132 314628
rect 394608 313216 394660 313268
rect 580816 313216 580868 313268
rect 393964 311856 394016 311908
rect 580172 311856 580224 311908
rect 32404 307708 32456 307760
rect 189080 307708 189132 307760
rect 394240 306280 394292 306332
rect 403624 306280 403676 306332
rect 3792 300772 3844 300824
rect 189080 300772 189132 300824
rect 394608 300772 394660 300824
rect 549904 300772 549956 300824
rect 3884 293904 3936 293956
rect 189080 293904 189132 293956
rect 394608 293904 394660 293956
rect 580908 293904 580960 293956
rect 394608 288328 394660 288380
rect 407764 288328 407816 288380
rect 3976 286968 4028 287020
rect 189080 286968 189132 287020
rect 393688 281256 393740 281308
rect 396724 281256 396776 281308
rect 17224 280100 17276 280152
rect 189080 280100 189132 280152
rect 394608 275952 394660 276004
rect 580264 275952 580316 276004
rect 10324 274592 10376 274644
rect 189080 274592 189132 274644
rect 3424 267656 3476 267708
rect 189080 267656 189132 267708
rect 394608 263508 394660 263560
rect 580356 263508 580408 263560
rect 3516 260788 3568 260840
rect 189080 260788 189132 260840
rect 394056 258068 394108 258120
rect 580172 258068 580224 258120
rect 394608 256640 394660 256692
rect 580448 256640 580500 256692
rect 4068 253852 4120 253904
rect 189080 253852 189132 253904
rect 3608 246984 3660 247036
rect 189080 246984 189132 247036
rect 394608 244196 394660 244248
rect 580540 244196 580592 244248
rect 3700 240048 3752 240100
rect 189080 240048 189132 240100
rect 394608 238688 394660 238740
rect 580264 238688 580316 238740
rect 3792 234540 3844 234592
rect 189080 234540 189132 234592
rect 393964 231820 394016 231872
rect 579804 231820 579856 231872
rect 3884 227672 3936 227724
rect 189080 227672 189132 227724
rect 394608 226244 394660 226296
rect 580356 226244 580408 226296
rect 3424 220736 3476 220788
rect 189080 220736 189132 220788
rect 393964 218016 394016 218068
rect 580172 218016 580224 218068
rect 3516 213868 3568 213920
rect 189080 213868 189132 213920
rect 3424 206932 3476 206984
rect 189080 206932 189132 206984
rect 394608 206252 394660 206304
rect 580172 206252 580224 206304
rect 3148 200064 3200 200116
rect 189080 200064 189132 200116
rect 3424 193196 3476 193248
rect 189080 193196 189132 193248
rect 394056 193128 394108 193180
rect 580172 193128 580224 193180
rect 3424 179392 3476 179444
rect 189080 179392 189132 179444
rect 393964 179324 394016 179376
rect 580172 179324 580224 179376
rect 394240 166948 394292 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 189816 164160 189868 164212
rect 3608 158720 3660 158772
rect 189080 158720 189132 158772
rect 394148 153144 394200 153196
rect 580172 153144 580224 153196
rect 3516 139408 3568 139460
rect 189080 139408 189132 139460
rect 394056 139340 394108 139392
rect 580172 139340 580224 139392
rect 3424 137912 3476 137964
rect 189724 137912 189776 137964
rect 393780 131112 393832 131164
rect 395344 131112 395396 131164
rect 393964 126896 394016 126948
rect 580172 126896 580224 126948
rect 3424 118668 3476 118720
rect 189080 118668 189132 118720
rect 395344 115200 395396 115252
rect 580264 115200 580316 115252
rect 394516 113092 394568 113144
rect 580172 113092 580224 113144
rect 394608 111800 394660 111852
rect 395344 111800 395396 111852
rect 3332 111732 3384 111784
rect 190184 111732 190236 111784
rect 224960 110168 225012 110220
rect 225144 110168 225196 110220
rect 238760 110168 238812 110220
rect 238944 110168 238996 110220
rect 345020 110168 345072 110220
rect 345204 110168 345256 110220
rect 285680 108808 285732 108860
rect 286324 108808 286376 108860
rect 314660 108808 314712 108860
rect 314844 108808 314896 108860
rect 390560 108672 390612 108724
rect 400864 108672 400916 108724
rect 188344 108604 188396 108656
rect 209596 108604 209648 108656
rect 339408 108604 339460 108656
rect 124220 108536 124272 108588
rect 234804 108536 234856 108588
rect 253204 108536 253256 108588
rect 262312 108536 262364 108588
rect 285956 108536 286008 108588
rect 290372 108536 290424 108588
rect 313096 108536 313148 108588
rect 117320 108468 117372 108520
rect 232320 108468 232372 108520
rect 235356 108468 235408 108520
rect 249800 108468 249852 108520
rect 250444 108468 250496 108520
rect 264336 108468 264388 108520
rect 278780 108468 278832 108520
rect 287888 108468 287940 108520
rect 110420 108400 110472 108452
rect 229928 108400 229980 108452
rect 247684 108400 247736 108452
rect 263140 108400 263192 108452
rect 265624 108400 265676 108452
rect 273812 108400 273864 108452
rect 273904 108400 273956 108452
rect 280160 108400 280212 108452
rect 281540 108400 281592 108452
rect 288716 108400 288768 108452
rect 302884 108400 302936 108452
rect 315304 108400 315356 108452
rect 333336 108400 333388 108452
rect 338672 108400 338724 108452
rect 17224 108332 17276 108384
rect 197452 108332 197504 108384
rect 235264 108332 235316 108384
rect 266820 108332 266872 108384
rect 277768 108332 277820 108384
rect 287520 108332 287572 108384
rect 300032 108332 300084 108384
rect 309784 108332 309836 108384
rect 310612 108332 310664 108384
rect 333244 108332 333296 108384
rect 10324 108264 10376 108316
rect 194232 108264 194284 108316
rect 218704 108264 218756 108316
rect 222200 108264 222252 108316
rect 223580 108264 223632 108316
rect 268844 108264 268896 108316
rect 274640 108264 274692 108316
rect 285680 108264 285732 108316
rect 304908 108264 304960 108316
rect 328460 108264 328512 108316
rect 381176 108604 381228 108656
rect 396724 108604 396776 108656
rect 370228 108536 370280 108588
rect 392584 108536 392636 108588
rect 429200 108468 429252 108520
rect 341892 108400 341944 108452
rect 436100 108400 436152 108452
rect 344284 108332 344336 108384
rect 443000 108332 443052 108384
rect 247224 108128 247276 108180
rect 248512 108128 248564 108180
rect 257436 108128 257488 108180
rect 258264 108128 258316 108180
rect 296720 108128 296772 108180
rect 297364 108128 297416 108180
rect 257344 108060 257396 108112
rect 259092 108060 259144 108112
rect 330116 108060 330168 108112
rect 337384 108060 337436 108112
rect 346768 108264 346820 108316
rect 449900 108264 449952 108316
rect 347044 108060 347096 108112
rect 252008 107992 252060 108044
rect 259552 107992 259604 108044
rect 295248 107992 295300 108044
rect 297364 107992 297416 108044
rect 319996 107924 320048 107976
rect 327632 107924 327684 107976
rect 238116 107788 238168 107840
rect 241244 107788 241296 107840
rect 287428 107788 287480 107840
rect 290740 107788 290792 107840
rect 193864 107720 193916 107772
rect 194968 107720 195020 107772
rect 203524 107720 203576 107772
rect 205180 107720 205232 107772
rect 220084 107720 220136 107772
rect 226616 107720 226668 107772
rect 238024 107720 238076 107772
rect 240416 107720 240468 107772
rect 288440 107720 288492 107772
rect 291108 107720 291160 107772
rect 298468 107720 298520 107772
rect 302884 107720 302936 107772
rect 308588 107720 308640 107772
rect 311256 107720 311308 107772
rect 365812 107720 365864 107772
rect 369124 107720 369176 107772
rect 383660 107720 383712 107772
rect 385868 107720 385920 107772
rect 193956 107652 194008 107704
rect 194600 107652 194652 107704
rect 203708 107652 203760 107704
rect 204720 107652 204772 107704
rect 211804 107652 211856 107704
rect 212816 107652 212868 107704
rect 213184 107652 213236 107704
rect 214104 107652 214156 107704
rect 214656 107652 214708 107704
rect 216128 107652 216180 107704
rect 217324 107652 217376 107704
rect 218152 107652 218204 107704
rect 221556 107652 221608 107704
rect 223028 107652 223080 107704
rect 235448 107652 235500 107704
rect 236368 107652 236420 107704
rect 236644 107652 236696 107704
rect 238392 107652 238444 107704
rect 242164 107652 242216 107704
rect 244924 107652 244976 107704
rect 250536 107652 250588 107704
rect 253388 107652 253440 107704
rect 256056 107652 256108 107704
rect 257068 107652 257120 107704
rect 264244 107652 264296 107704
rect 265164 107652 265216 107704
rect 268384 107652 268436 107704
rect 269212 107652 269264 107704
rect 269764 107652 269816 107704
rect 270500 107652 270552 107704
rect 271144 107652 271196 107704
rect 272064 107652 272116 107704
rect 289084 107652 289136 107704
rect 289912 107652 289964 107704
rect 292396 107652 292448 107704
rect 292672 107652 292724 107704
rect 294788 107652 294840 107704
rect 295984 107652 296036 107704
rect 297272 107652 297324 107704
rect 300032 107652 300084 107704
rect 308220 107652 308272 107704
rect 309968 107652 310020 107704
rect 316684 107652 316736 107704
rect 319444 107652 319496 107704
rect 321560 107652 321612 107704
rect 323584 107652 323636 107704
rect 326436 107652 326488 107704
rect 327816 107652 327868 107704
rect 348332 107652 348384 107704
rect 351184 107652 351236 107704
rect 352012 107652 352064 107704
rect 353944 107652 353996 107704
rect 366640 107652 366692 107704
rect 367744 107652 367796 107704
rect 379980 107652 380032 107704
rect 381544 107652 381596 107704
rect 384028 107652 384080 107704
rect 385684 107652 385736 107704
rect 387340 107652 387392 107704
rect 392676 107652 392728 107704
rect 215392 107108 215444 107160
rect 215576 107108 215628 107160
rect 157340 107040 157392 107092
rect 246120 107040 246172 107092
rect 339868 107040 339920 107092
rect 430580 107040 430632 107092
rect 125600 106972 125652 107024
rect 234896 106972 234948 107024
rect 356888 106972 356940 107024
rect 480260 106972 480312 107024
rect 74540 106904 74592 106956
rect 217692 106904 217744 106956
rect 259460 106904 259512 106956
rect 281448 106904 281500 106956
rect 309416 106904 309468 106956
rect 340880 106904 340932 106956
rect 379612 106904 379664 106956
rect 546500 106904 546552 106956
rect 201500 106836 201552 106888
rect 202052 106836 202104 106888
rect 223764 106836 223816 106888
rect 224316 106836 224368 106888
rect 256884 106836 256936 106888
rect 257620 106836 257672 106888
rect 281724 106836 281776 106888
rect 282276 106836 282328 106888
rect 300860 106836 300912 106888
rect 301412 106836 301464 106888
rect 305092 106836 305144 106888
rect 305828 106836 305880 106888
rect 335360 106836 335412 106888
rect 335912 106836 335964 106888
rect 342260 106836 342312 106888
rect 342812 106836 342864 106888
rect 345112 106836 345164 106888
rect 346032 106836 346084 106888
rect 349344 106836 349396 106888
rect 349620 106836 349672 106888
rect 353392 106836 353444 106888
rect 354128 106836 354180 106888
rect 354772 106836 354824 106888
rect 355324 106836 355376 106888
rect 191840 106768 191892 106820
rect 192668 106768 192720 106820
rect 201592 106768 201644 106820
rect 202420 106768 202472 106820
rect 215392 106768 215444 106820
rect 216220 106768 216272 106820
rect 219440 106768 219492 106820
rect 220268 106768 220320 106820
rect 222292 106768 222344 106820
rect 223120 106768 223172 106820
rect 223672 106768 223724 106820
rect 223948 106768 224000 106820
rect 245752 106768 245804 106820
rect 246580 106768 246632 106820
rect 247132 106768 247184 106820
rect 247868 106768 247920 106820
rect 249892 106768 249944 106820
rect 250720 106768 250772 106820
rect 253940 106768 253992 106820
rect 254768 106768 254820 106820
rect 255320 106768 255372 106820
rect 255964 106768 256016 106820
rect 256792 106768 256844 106820
rect 257160 106768 257212 106820
rect 259552 106768 259604 106820
rect 260380 106768 260432 106820
rect 273352 106768 273404 106820
rect 274180 106768 274232 106820
rect 277584 106768 277636 106820
rect 278228 106768 278280 106820
rect 278872 106768 278924 106820
rect 279516 106768 279568 106820
rect 281632 106768 281684 106820
rect 281908 106768 281960 106820
rect 284392 106768 284444 106820
rect 285220 106768 285272 106820
rect 291200 106768 291252 106820
rect 291660 106768 291712 106820
rect 295432 106768 295484 106820
rect 296076 106768 296128 106820
rect 296812 106768 296864 106820
rect 297732 106768 297784 106820
rect 298100 106768 298152 106820
rect 299020 106768 299072 106820
rect 301044 106768 301096 106820
rect 301780 106768 301832 106820
rect 302240 106768 302292 106820
rect 303068 106768 303120 106820
rect 303712 106768 303764 106820
rect 304264 106768 304316 106820
rect 305000 106768 305052 106820
rect 305460 106768 305512 106820
rect 306380 106768 306432 106820
rect 307116 106768 307168 106820
rect 310520 106768 310572 106820
rect 311532 106768 311584 106820
rect 324320 106768 324372 106820
rect 325332 106768 325384 106820
rect 327172 106768 327224 106820
rect 327724 106768 327776 106820
rect 328552 106768 328604 106820
rect 329380 106768 329432 106820
rect 329840 106768 329892 106820
rect 330668 106768 330720 106820
rect 332600 106768 332652 106820
rect 333428 106768 333480 106820
rect 335544 106768 335596 106820
rect 336280 106768 336332 106820
rect 336740 106768 336792 106820
rect 337108 106768 337160 106820
rect 338212 106768 338264 106820
rect 338764 106768 338816 106820
rect 339500 106768 339552 106820
rect 340328 106768 340380 106820
rect 342444 106768 342496 106820
rect 343180 106768 343232 106820
rect 345204 106768 345256 106820
rect 345572 106768 345624 106820
rect 349160 106768 349212 106820
rect 350080 106768 350132 106820
rect 350540 106768 350592 106820
rect 351276 106768 351328 106820
rect 352012 106768 352064 106820
rect 352932 106768 352984 106820
rect 353300 106768 353352 106820
rect 353760 106768 353812 106820
rect 354680 106768 354732 106820
rect 354956 106768 355008 106820
rect 356060 106768 356112 106820
rect 356244 106768 356296 106820
rect 358820 106768 358872 106820
rect 359832 106768 359884 106820
rect 389272 106768 389324 106820
rect 389824 106768 389876 106820
rect 390560 106768 390612 106820
rect 391480 106768 391532 106820
rect 218244 106700 218296 106752
rect 219072 106700 219124 106752
rect 252744 106700 252796 106752
rect 253572 106700 253624 106752
rect 342352 106700 342404 106752
rect 342628 106700 342680 106752
rect 336832 106632 336884 106684
rect 337476 106632 337528 106684
rect 197452 106088 197504 106140
rect 198004 106088 198056 106140
rect 331220 106088 331272 106140
rect 331404 106088 331456 106140
rect 323032 105816 323084 105868
rect 323676 105816 323728 105868
rect 169760 105680 169812 105732
rect 250628 105680 250680 105732
rect 328920 105680 328972 105732
rect 398840 105680 398892 105732
rect 160100 105612 160152 105664
rect 247316 105612 247368 105664
rect 358084 105612 358136 105664
rect 483020 105612 483072 105664
rect 60740 105544 60792 105596
rect 212908 105544 212960 105596
rect 324412 105544 324464 105596
rect 324596 105544 324648 105596
rect 380440 105544 380492 105596
rect 547880 105544 547932 105596
rect 363236 105408 363288 105460
rect 363512 105408 363564 105460
rect 351920 104728 351972 104780
rect 352564 104728 352616 104780
rect 243084 104592 243136 104644
rect 382372 104592 382424 104644
rect 386604 104592 386656 104644
rect 252560 104456 252612 104508
rect 252836 104456 252888 104508
rect 317512 104456 317564 104508
rect 317696 104456 317748 104508
rect 378140 104456 378192 104508
rect 378416 104456 378468 104508
rect 243084 104388 243136 104440
rect 382372 104388 382424 104440
rect 386604 104388 386656 104440
rect 211436 104320 211488 104372
rect 211620 104320 211672 104372
rect 263876 104320 263928 104372
rect 264060 104320 264112 104372
rect 317420 104320 317472 104372
rect 317604 104320 317656 104372
rect 385132 104320 385184 104372
rect 385776 104320 385828 104372
rect 173900 104252 173952 104304
rect 251824 104252 251876 104304
rect 331312 104252 331364 104304
rect 405740 104252 405792 104304
rect 164240 104184 164292 104236
rect 247224 104184 247276 104236
rect 263692 104184 263744 104236
rect 264428 104184 264480 104236
rect 265072 104184 265124 104236
rect 265716 104184 265768 104236
rect 266544 104184 266596 104236
rect 267372 104184 267424 104236
rect 270684 104184 270736 104236
rect 271420 104184 271472 104236
rect 271972 104184 272024 104236
rect 272616 104184 272668 104236
rect 277400 104184 277452 104236
rect 277860 104184 277912 104236
rect 313372 104184 313424 104236
rect 313924 104184 313976 104236
rect 314660 104184 314712 104236
rect 315212 104184 315264 104236
rect 317420 104184 317472 104236
rect 318064 104184 318116 104236
rect 359280 104184 359332 104236
rect 487160 104184 487212 104236
rect 57980 104116 58032 104168
rect 205640 104048 205692 104100
rect 206468 104048 206520 104100
rect 207020 104116 207072 104168
rect 207664 104116 207716 104168
rect 209780 104116 209832 104168
rect 210516 104116 210568 104168
rect 211252 104116 211304 104168
rect 212172 104116 212224 104168
rect 214012 104116 214064 104168
rect 214564 104116 214616 104168
rect 225052 104116 225104 104168
rect 225604 104116 225656 104168
rect 227720 104116 227772 104168
rect 228364 104116 228416 104168
rect 229284 104116 229336 104168
rect 230020 104116 230072 104168
rect 232044 104116 232096 104168
rect 232412 104116 232464 104168
rect 233332 104116 233384 104168
rect 234068 104116 234120 104168
rect 238852 104116 238904 104168
rect 239312 104116 239364 104168
rect 242992 104116 243044 104168
rect 243820 104116 243872 104168
rect 247040 104116 247092 104168
rect 276940 104116 276992 104168
rect 363052 104116 363104 104168
rect 363420 104116 363472 104168
rect 364340 104116 364392 104168
rect 364708 104116 364760 104168
rect 367100 104116 367152 104168
rect 367560 104116 367612 104168
rect 369860 104116 369912 104168
rect 370780 104116 370832 104168
rect 371240 104116 371292 104168
rect 371976 104116 372028 104168
rect 372620 104116 372672 104168
rect 373632 104116 373684 104168
rect 374000 104116 374052 104168
rect 374828 104116 374880 104168
rect 376760 104116 376812 104168
rect 377220 104116 377272 104168
rect 378232 104116 378284 104168
rect 378876 104116 378928 104168
rect 212080 104048 212132 104100
rect 231952 104048 232004 104100
rect 232780 104048 232832 104100
rect 362960 104048 363012 104100
rect 363880 104048 363932 104100
rect 364432 104048 364484 104100
rect 365076 104048 365128 104100
rect 377128 104048 377180 104100
rect 539600 104116 539652 104168
rect 385040 104048 385092 104100
rect 385408 104048 385460 104100
rect 386512 104048 386564 104100
rect 387432 104048 387484 104100
rect 387984 104048 388036 104100
rect 388628 104048 388680 104100
rect 299480 103912 299532 103964
rect 300124 103912 300176 103964
rect 276020 103504 276072 103556
rect 276204 103504 276256 103556
rect 187700 102892 187752 102944
rect 256976 102892 257028 102944
rect 171140 102824 171192 102876
rect 249892 102824 249944 102876
rect 349436 102824 349488 102876
rect 458180 102824 458232 102876
rect 46940 102756 46992 102808
rect 208308 102756 208360 102808
rect 360292 102756 360344 102808
rect 489920 102756 489972 102808
rect 361580 102144 361632 102196
rect 362316 102144 362368 102196
rect 175280 101532 175332 101584
rect 251364 101532 251416 101584
rect 131120 101464 131172 101516
rect 236920 101464 236972 101516
rect 361764 101464 361816 101516
rect 494060 101464 494112 101516
rect 14464 101396 14516 101448
rect 194692 101396 194744 101448
rect 225144 101396 225196 101448
rect 225972 101396 226024 101448
rect 230388 101396 230440 101448
rect 230572 101396 230624 101448
rect 242900 101396 242952 101448
rect 243176 101396 243228 101448
rect 251180 101396 251232 101448
rect 277400 101396 277452 101448
rect 315580 101396 315632 101448
rect 360292 101396 360344 101448
rect 368480 101396 368532 101448
rect 368664 101396 368716 101448
rect 375472 101396 375524 101448
rect 534080 101396 534132 101448
rect 382280 101328 382332 101380
rect 382464 101328 382516 101380
rect 229192 100920 229244 100972
rect 229468 100920 229520 100972
rect 238944 100716 238996 100768
rect 239772 100716 239824 100768
rect 394424 100648 394476 100700
rect 580172 100648 580224 100700
rect 178040 100104 178092 100156
rect 250536 100104 250588 100156
rect 151820 100036 151872 100088
rect 244372 100036 244424 100088
rect 327264 100036 327316 100088
rect 394700 100036 394752 100088
rect 29000 99968 29052 100020
rect 201500 99968 201552 100020
rect 347872 99968 347924 100020
rect 456892 99968 456944 100020
rect 386420 99696 386472 99748
rect 386696 99696 386748 99748
rect 236092 99220 236144 99272
rect 236460 99220 236512 99272
rect 182180 98744 182232 98796
rect 254124 98744 254176 98796
rect 329932 98744 329984 98796
rect 402980 98744 403032 98796
rect 81440 98676 81492 98728
rect 219624 98676 219676 98728
rect 363512 98676 363564 98728
rect 498200 98676 498252 98728
rect 6920 98608 6972 98660
rect 193956 98608 194008 98660
rect 382464 98608 382516 98660
rect 556160 98608 556212 98660
rect 184940 97384 184992 97436
rect 255504 97384 255556 97436
rect 142160 97316 142212 97368
rect 240232 97316 240284 97368
rect 343640 97316 343692 97368
rect 441620 97316 441672 97368
rect 8300 97248 8352 97300
rect 193864 97248 193916 97300
rect 367744 97248 367796 97300
rect 507860 97248 507912 97300
rect 193404 96024 193456 96076
rect 257436 96024 257488 96076
rect 328736 96024 328788 96076
rect 398932 96024 398984 96076
rect 129740 95956 129792 96008
rect 236092 95956 236144 96008
rect 336924 95956 336976 96008
rect 422300 95956 422352 96008
rect 34520 95888 34572 95940
rect 203064 95888 203116 95940
rect 375472 95888 375524 95940
rect 536840 95888 536892 95940
rect 128360 94528 128412 94580
rect 235448 94528 235500 94580
rect 352104 94528 352156 94580
rect 466460 94528 466512 94580
rect 78680 94460 78732 94512
rect 218244 94460 218296 94512
rect 321744 94460 321796 94512
rect 380992 94460 381044 94512
rect 381544 94460 381596 94512
rect 547972 94460 548024 94512
rect 325792 93236 325844 93288
rect 391940 93236 391992 93288
rect 132500 93168 132552 93220
rect 237472 93168 237524 93220
rect 335636 93168 335688 93220
rect 418160 93168 418212 93220
rect 89720 93100 89772 93152
rect 221464 93100 221516 93152
rect 385776 93100 385828 93152
rect 557540 93100 557592 93152
rect 135260 91808 135312 91860
rect 239036 91808 239088 91860
rect 341156 91808 341208 91860
rect 434720 91808 434772 91860
rect 35900 91740 35952 91792
rect 203616 91740 203668 91792
rect 307852 91740 307904 91792
rect 340972 91740 341024 91792
rect 383752 91740 383804 91792
rect 561680 91740 561732 91792
rect 139400 90380 139452 90432
rect 238944 90380 238996 90432
rect 350724 90380 350776 90432
rect 463700 90380 463752 90432
rect 48320 90312 48372 90364
rect 208492 90312 208544 90364
rect 316132 90312 316184 90364
rect 364524 90312 364576 90364
rect 385132 90312 385184 90364
rect 564440 90312 564492 90364
rect 143540 89020 143592 89072
rect 238116 89020 238168 89072
rect 329840 89020 329892 89072
rect 404360 89020 404412 89072
rect 62120 88952 62172 89004
rect 212724 88952 212776 89004
rect 324596 88952 324648 89004
rect 387800 88952 387852 89004
rect 388076 88952 388128 89004
rect 571984 88952 572036 89004
rect 146300 87660 146352 87712
rect 241704 87660 241756 87712
rect 345296 87660 345348 87712
rect 445760 87660 445812 87712
rect 77300 87592 77352 87644
rect 218152 87592 218204 87644
rect 389364 87592 389416 87644
rect 575480 87592 575532 87644
rect 394332 86912 394384 86964
rect 580172 86912 580224 86964
rect 150440 86300 150492 86352
rect 243176 86300 243228 86352
rect 114560 86232 114612 86284
rect 230664 86232 230716 86284
rect 327172 86232 327224 86284
rect 396080 86232 396132 86284
rect 3332 85484 3384 85536
rect 190092 85484 190144 85536
rect 179420 84872 179472 84924
rect 252744 84872 252796 84924
rect 337384 84872 337436 84924
rect 401600 84872 401652 84924
rect 92480 84804 92532 84856
rect 223856 84804 223908 84856
rect 361672 84804 361724 84856
rect 495440 84804 495492 84856
rect 153200 83512 153252 83564
rect 242164 83512 242216 83564
rect 331404 83512 331456 83564
rect 408500 83512 408552 83564
rect 102140 83444 102192 83496
rect 226432 83444 226484 83496
rect 369124 83444 369176 83496
rect 506480 83444 506532 83496
rect 126980 82152 127032 82204
rect 234712 82152 234764 82204
rect 334164 82152 334216 82204
rect 415400 82152 415452 82204
rect 56600 82084 56652 82136
rect 211344 82084 211396 82136
rect 365812 82084 365864 82136
rect 509240 82084 509292 82136
rect 161480 80724 161532 80776
rect 247224 80724 247276 80776
rect 338304 80724 338356 80776
rect 426440 80724 426492 80776
rect 66260 80656 66312 80708
rect 214012 80656 214064 80708
rect 370044 80656 370096 80708
rect 520280 80656 520332 80708
rect 165620 79364 165672 79416
rect 248512 79364 248564 79416
rect 342536 79364 342588 79416
rect 437480 79364 437532 79416
rect 18604 79296 18656 79348
rect 197544 79296 197596 79348
rect 369952 79296 370004 79348
rect 517520 79296 517572 79348
rect 254124 78140 254176 78192
rect 279056 78140 279108 78192
rect 183560 78004 183612 78056
rect 253940 78004 253992 78056
rect 342444 78004 342496 78056
rect 440332 78004 440384 78056
rect 75920 77936 75972 77988
rect 217324 77936 217376 77988
rect 369860 77936 369912 77988
rect 521660 77936 521712 77988
rect 133880 76576 133932 76628
rect 237564 76576 237616 76628
rect 343732 76576 343784 76628
rect 444380 76576 444432 76628
rect 63500 76508 63552 76560
rect 213184 76508 213236 76560
rect 309232 76508 309284 76560
rect 343640 76508 343692 76560
rect 372896 76508 372948 76560
rect 528560 76508 528612 76560
rect 147680 75216 147732 75268
rect 243084 75216 243136 75268
rect 345204 75216 345256 75268
rect 448520 75216 448572 75268
rect 52460 75148 52512 75200
rect 209964 75148 210016 75200
rect 375380 75148 375432 75200
rect 535460 75148 535512 75200
rect 151912 73856 151964 73908
rect 242992 73856 243044 73908
rect 351184 73856 351236 73908
rect 455420 73856 455472 73908
rect 49700 73788 49752 73840
rect 208584 73788 208636 73840
rect 311992 73788 312044 73840
rect 350724 73788 350776 73840
rect 378324 73788 378376 73840
rect 542360 73788 542412 73840
rect 394240 73108 394292 73160
rect 579988 73108 580040 73160
rect 154580 72496 154632 72548
rect 244464 72496 244516 72548
rect 44180 72428 44232 72480
rect 207204 72428 207256 72480
rect 323124 72428 323176 72480
rect 382464 72428 382516 72480
rect 3332 71680 3384 71732
rect 190000 71680 190052 71732
rect 353944 71068 353996 71120
rect 465172 71068 465224 71120
rect 185032 71000 185084 71052
rect 255412 71000 255464 71052
rect 379520 71000 379572 71052
rect 549260 71000 549312 71052
rect 162860 69708 162912 69760
rect 247132 69708 247184 69760
rect 352012 69708 352064 69760
rect 469220 69708 469272 69760
rect 41420 69640 41472 69692
rect 205824 69640 205876 69692
rect 381084 69640 381136 69692
rect 553400 69640 553452 69692
rect 167000 68348 167052 68400
rect 248604 68348 248656 68400
rect 356244 68348 356296 68400
rect 481640 68348 481692 68400
rect 27620 68280 27672 68332
rect 201684 68280 201736 68332
rect 383660 68280 383712 68332
rect 560300 68280 560352 68332
rect 180800 66920 180852 66972
rect 254032 66920 254084 66972
rect 91100 66852 91152 66904
rect 222292 66852 222344 66904
rect 314844 66852 314896 66904
rect 357440 66852 357492 66904
rect 357624 66852 357676 66904
rect 484400 66852 484452 66904
rect 135352 65560 135404 65612
rect 236644 65560 236696 65612
rect 95240 65492 95292 65544
rect 225236 65492 225288 65544
rect 359004 65492 359056 65544
rect 488540 65492 488592 65544
rect 138020 64200 138072 64252
rect 238852 64200 238904 64252
rect 99380 64132 99432 64184
rect 225144 64132 225196 64184
rect 363144 64132 363196 64184
rect 498292 64132 498344 64184
rect 155960 62840 156012 62892
rect 245844 62840 245896 62892
rect 331312 62840 331364 62892
rect 407120 62840 407172 62892
rect 21364 62772 21416 62824
rect 196164 62772 196216 62824
rect 364616 62772 364668 62824
rect 502340 62772 502392 62824
rect 69020 61344 69072 61396
rect 215484 61344 215536 61396
rect 310704 61344 310756 61396
rect 347872 61344 347924 61396
rect 367284 61344 367336 61396
rect 513380 61344 513432 61396
rect 394148 60664 394200 60716
rect 580172 60664 580224 60716
rect 71780 59984 71832 60036
rect 216772 59984 216824 60036
rect 328644 59984 328696 60036
rect 397460 59984 397512 60036
rect 85580 58624 85632 58676
rect 221004 58624 221056 58676
rect 317696 58624 317748 58676
rect 368664 58624 368716 58676
rect 368756 58624 368808 58676
rect 516140 58624 516192 58676
rect 328552 57264 328604 57316
rect 400220 57264 400272 57316
rect 100760 57196 100812 57248
rect 220084 57196 220136 57248
rect 385684 57196 385736 57248
rect 558920 57196 558972 57248
rect 110512 55836 110564 55888
rect 229284 55836 229336 55888
rect 324504 55836 324556 55888
rect 385132 55836 385184 55888
rect 385224 55836 385276 55888
rect 563060 55836 563112 55888
rect 160192 54544 160244 54596
rect 245752 54544 245804 54596
rect 324412 54544 324464 54596
rect 386696 54544 386748 54596
rect 88340 54476 88392 54528
rect 222384 54476 222436 54528
rect 386604 54476 386656 54528
rect 565820 54476 565872 54528
rect 149060 53116 149112 53168
rect 242900 53116 242952 53168
rect 102232 53048 102284 53100
rect 226524 53048 226576 53100
rect 321652 53048 321704 53100
rect 379520 53048 379572 53100
rect 386512 53048 386564 53100
rect 569960 53048 570012 53100
rect 219624 51756 219676 51808
rect 266544 51756 266596 51808
rect 121460 51688 121512 51740
rect 233424 51688 233476 51740
rect 320364 51688 320416 51740
rect 375380 51688 375432 51740
rect 387984 51688 388036 51740
rect 572076 51688 572128 51740
rect 144920 50328 144972 50380
rect 241612 50328 241664 50380
rect 317604 50328 317656 50380
rect 365812 50328 365864 50380
rect 389272 50328 389324 50380
rect 574744 50328 574796 50380
rect 346492 49036 346544 49088
rect 452660 49036 452712 49088
rect 59360 48968 59412 49020
rect 211252 48968 211304 49020
rect 216772 48968 216824 49020
rect 266452 48968 266504 49020
rect 389180 48968 389232 49020
rect 574100 48968 574152 49020
rect 209964 47608 210016 47660
rect 263784 47608 263836 47660
rect 349344 47608 349396 47660
rect 459560 47608 459612 47660
rect 86960 47540 87012 47592
rect 218704 47540 218756 47592
rect 400864 47540 400916 47592
rect 578240 47540 578292 47592
rect 143632 46180 143684 46232
rect 241520 46180 241572 46232
rect 353484 46180 353536 46232
rect 470600 46180 470652 46232
rect 3516 45500 3568 45552
rect 189908 45500 189960 45552
rect 205824 44820 205876 44872
rect 262312 44820 262364 44872
rect 356152 44820 356204 44872
rect 477500 44820 477552 44872
rect 199016 43460 199068 43512
rect 259736 43460 259788 43512
rect 30380 43392 30432 43444
rect 201592 43392 201644 43444
rect 357532 43392 357584 43444
rect 481732 43392 481784 43444
rect 176660 42100 176712 42152
rect 252652 42100 252704 42152
rect 70400 42032 70452 42084
rect 215392 42032 215444 42084
rect 358912 42032 358964 42084
rect 485780 42032 485832 42084
rect 158720 40672 158772 40724
rect 245936 40672 245988 40724
rect 363052 40672 363104 40724
rect 499580 40672 499632 40724
rect 127072 39312 127124 39364
rect 236276 39312 236328 39364
rect 242900 39312 242952 39364
rect 274916 39312 274968 39364
rect 365720 39312 365772 39364
rect 506572 39312 506624 39364
rect 136640 37884 136692 37936
rect 238760 37884 238812 37936
rect 316040 37884 316092 37936
rect 361672 37884 361724 37936
rect 368572 37884 368624 37936
rect 514760 37884 514812 37936
rect 236000 36592 236052 36644
rect 273444 36592 273496 36644
rect 140780 36524 140832 36576
rect 238024 36524 238076 36576
rect 314752 36524 314804 36576
rect 357532 36524 357584 36576
rect 361580 36524 361632 36576
rect 496820 36524 496872 36576
rect 118700 35164 118752 35216
rect 232044 35164 232096 35216
rect 233424 35164 233476 35216
rect 271144 35164 271196 35216
rect 313464 35164 313516 35216
rect 354956 35164 355008 35216
rect 358820 35164 358872 35216
rect 490012 35164 490064 35216
rect 345112 33804 345164 33856
rect 448612 33804 448664 33856
rect 17960 33736 18012 33788
rect 197452 33736 197504 33788
rect 197544 33736 197596 33788
rect 259644 33736 259696 33788
rect 386420 33736 386472 33788
rect 567200 33736 567252 33788
rect 2872 33056 2924 33108
rect 189816 33056 189868 33108
rect 394056 33056 394108 33108
rect 580172 33056 580224 33108
rect 189080 32376 189132 32428
rect 255964 32376 256016 32428
rect 324320 32376 324372 32428
rect 389180 32376 389232 32428
rect 215392 31084 215444 31136
rect 265072 31084 265124 31136
rect 73160 31016 73212 31068
rect 216864 31016 216916 31068
rect 307760 31016 307812 31068
rect 336924 31016 336976 31068
rect 371424 31016 371476 31068
rect 523040 31016 523092 31068
rect 193496 29656 193548 29708
rect 258172 29656 258224 29708
rect 338764 29656 338816 29708
rect 411260 29656 411312 29708
rect 60832 29588 60884 29640
rect 211804 29588 211856 29640
rect 311900 29588 311952 29640
rect 349344 29588 349396 29640
rect 395344 29588 395396 29640
rect 580264 29588 580316 29640
rect 310612 28432 310664 28484
rect 346492 28432 346544 28484
rect 190460 28296 190512 28348
rect 256792 28296 256844 28348
rect 346400 28296 346452 28348
rect 451280 28296 451332 28348
rect 67640 28228 67692 28280
rect 215576 28228 215628 28280
rect 387892 28228 387944 28280
rect 570604 28228 570656 28280
rect 186320 26936 186372 26988
rect 255320 26936 255372 26988
rect 341064 26936 341116 26988
rect 433340 26936 433392 26988
rect 77392 26868 77444 26920
rect 218336 26868 218388 26920
rect 305184 26868 305236 26920
rect 329840 26868 329892 26920
rect 385040 26868 385092 26920
rect 564532 26868 564584 26920
rect 176752 25576 176804 25628
rect 252836 25576 252888 25628
rect 311164 25576 311216 25628
rect 339684 25576 339736 25628
rect 85672 25508 85724 25560
rect 220912 25508 220964 25560
rect 258080 25508 258132 25560
rect 280252 25508 280304 25560
rect 325700 25508 325752 25560
rect 390836 25508 390888 25560
rect 392676 25508 392728 25560
rect 568580 25508 568632 25560
rect 323032 24148 323084 24200
rect 383660 24148 383712 24200
rect 172520 24080 172572 24132
rect 251272 24080 251324 24132
rect 261116 24080 261168 24132
rect 281816 24080 281868 24132
rect 382372 24080 382424 24132
rect 554780 24080 554832 24132
rect 314660 22788 314712 22840
rect 358820 22788 358872 22840
rect 168380 22720 168432 22772
rect 249984 22720 250036 22772
rect 252560 22720 252612 22772
rect 278964 22720 279016 22772
rect 298192 22720 298244 22772
rect 310612 22720 310664 22772
rect 327080 22720 327132 22772
rect 393320 22720 393372 22772
rect 396724 22720 396776 22772
rect 550640 22720 550692 22772
rect 302332 21564 302384 21616
rect 321652 21564 321704 21616
rect 321560 21428 321612 21480
rect 378324 21428 378376 21480
rect 55220 21360 55272 21412
rect 211436 21360 211488 21412
rect 214012 21360 214064 21412
rect 265164 21360 265216 21412
rect 371332 21360 371384 21412
rect 523132 21360 523184 21412
rect 393964 20612 394016 20664
rect 580172 20612 580224 20664
rect 210056 20000 210108 20052
rect 250444 20000 250496 20052
rect 319444 20000 319496 20052
rect 363052 20000 363104 20052
rect 192116 19932 192168 19984
rect 256884 19932 256936 19984
rect 334072 19932 334124 19984
rect 415492 19932 415544 19984
rect 203064 18640 203116 18692
rect 261024 18640 261076 18692
rect 309876 18640 309928 18692
rect 338304 18640 338356 18692
rect 69112 18572 69164 18624
rect 214564 18572 214616 18624
rect 263784 18572 263836 18624
rect 281724 18572 281776 18624
rect 327816 18572 327868 18624
rect 390928 18572 390980 18624
rect 392584 18572 392636 18624
rect 518900 18572 518952 18624
rect 200396 17280 200448 17332
rect 259552 17280 259604 17332
rect 315304 17280 315356 17332
rect 323032 17280 323084 17332
rect 323584 17280 323636 17332
rect 377036 17280 377088 17332
rect 37280 17212 37332 17264
rect 203524 17212 203576 17264
rect 218060 17212 218112 17264
rect 266636 17212 266688 17264
rect 301136 17212 301188 17264
rect 317604 17212 317656 17264
rect 362960 17212 363012 17264
rect 500960 17212 501012 17264
rect 211712 15920 211764 15972
rect 263692 15920 263744 15972
rect 303804 15920 303856 15972
rect 326344 15920 326396 15972
rect 51080 15852 51132 15904
rect 188344 15852 188396 15904
rect 196808 15852 196860 15904
rect 251824 15852 251876 15904
rect 256700 15852 256752 15904
rect 273904 15852 273956 15904
rect 313372 15852 313424 15904
rect 356336 15852 356388 15904
rect 368480 15852 368532 15904
rect 515496 15852 515548 15904
rect 306472 14560 306524 14612
rect 333888 14560 333940 14612
rect 221096 14492 221148 14544
rect 267832 14492 267884 14544
rect 327724 14492 327776 14544
rect 372896 14492 372948 14544
rect 168472 14424 168524 14476
rect 235356 14424 235408 14476
rect 306564 14424 306616 14476
rect 334624 14424 334676 14476
rect 364432 14424 364484 14476
rect 505376 14424 505428 14476
rect 123024 13336 123076 13388
rect 233332 13336 233384 13388
rect 119896 13268 119948 13320
rect 231952 13268 232004 13320
rect 116400 13200 116452 13252
rect 232136 13200 232188 13252
rect 367192 13200 367244 13252
rect 511264 13200 511316 13252
rect 112352 13132 112404 13184
rect 230572 13132 230624 13184
rect 303712 13132 303764 13184
rect 328000 13132 328052 13184
rect 371240 13132 371292 13184
rect 525432 13132 525484 13184
rect 22560 13064 22612 13116
rect 198924 13064 198976 13116
rect 232044 13064 232096 13116
rect 270684 13064 270736 13116
rect 270776 13064 270828 13116
rect 284576 13064 284628 13116
rect 317512 13064 317564 13116
rect 365720 13064 365772 13116
rect 374184 13064 374236 13116
rect 532056 13064 532108 13116
rect 109040 12044 109092 12096
rect 229192 12044 229244 12096
rect 105728 11976 105780 12028
rect 227904 11976 227956 12028
rect 98184 11908 98236 11960
rect 225052 11908 225104 11960
rect 93860 11840 93912 11892
rect 223764 11840 223816 11892
rect 354864 11840 354916 11892
rect 474096 11840 474148 11892
rect 84200 11772 84252 11824
rect 220820 11772 220872 11824
rect 240140 11772 240192 11824
rect 273352 11772 273404 11824
rect 301044 11772 301096 11824
rect 320456 11772 320508 11824
rect 360384 11772 360436 11824
rect 493048 11772 493100 11824
rect 80888 11704 80940 11756
rect 219532 11704 219584 11756
rect 228272 11704 228324 11756
rect 269764 11704 269816 11756
rect 310520 11704 310572 11756
rect 349344 11704 349396 11756
rect 364340 11704 364392 11756
rect 503720 11704 503772 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 168380 11636 168432 11688
rect 169576 11636 169628 11688
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 331220 10820 331272 10872
rect 407212 10820 407264 10872
rect 332692 10752 332744 10804
rect 410800 10752 410852 10804
rect 333980 10684 334032 10736
rect 414296 10684 414348 10736
rect 108120 10616 108172 10668
rect 229376 10616 229428 10668
rect 335452 10616 335504 10668
rect 417424 10616 417476 10668
rect 104072 10548 104124 10600
rect 227812 10548 227864 10600
rect 335544 10548 335596 10600
rect 420920 10548 420972 10600
rect 97448 10480 97500 10532
rect 224960 10480 225012 10532
rect 336832 10480 336884 10532
rect 423680 10480 423732 10532
rect 93952 10412 94004 10464
rect 223672 10412 223724 10464
rect 267740 10412 267792 10464
rect 283104 10412 283156 10464
rect 338212 10412 338264 10464
rect 428464 10412 428516 10464
rect 52552 10344 52604 10396
rect 209872 10344 209924 10396
rect 226340 10344 226392 10396
rect 269212 10344 269264 10396
rect 302240 10344 302292 10396
rect 324412 10344 324464 10396
rect 339592 10344 339644 10396
rect 432052 10344 432104 10396
rect 44272 10276 44324 10328
rect 207112 10276 207164 10328
rect 225144 10276 225196 10328
rect 268384 10276 268436 10328
rect 305092 10276 305144 10328
rect 332692 10276 332744 10328
rect 342352 10276 342404 10328
rect 439136 10276 439188 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 309784 9596 309836 9648
rect 315028 9596 315080 9648
rect 322940 9392 322992 9444
rect 382372 9392 382424 9444
rect 372804 9324 372856 9376
rect 527824 9324 527876 9376
rect 374092 9256 374144 9308
rect 531320 9256 531372 9308
rect 376852 9188 376904 9240
rect 538404 9188 538456 9240
rect 376944 9120 376996 9172
rect 541992 9120 542044 9172
rect 239312 9052 239364 9104
rect 265624 9052 265676 9104
rect 317420 9052 317472 9104
rect 368204 9052 368256 9104
rect 378232 9052 378284 9104
rect 545488 9052 545540 9104
rect 40684 8984 40736 9036
rect 205732 8984 205784 9036
rect 208584 8984 208636 9036
rect 263876 8984 263928 9036
rect 302884 8984 302936 9036
rect 13544 8916 13596 8968
rect 196072 8916 196124 8968
rect 202696 8916 202748 8968
rect 260932 8916 260984 8968
rect 295524 8916 295576 8968
rect 303160 8916 303212 8968
rect 318892 8984 318944 9036
rect 371700 8984 371752 9036
rect 380900 8984 380952 9036
rect 552664 8984 552716 9036
rect 310244 8916 310296 8968
rect 320272 8916 320324 8968
rect 375288 8916 375340 8968
rect 382280 8916 382332 8968
rect 556160 8916 556212 8968
rect 83280 7828 83332 7880
rect 219440 7828 219492 7880
rect 33600 7760 33652 7812
rect 202972 7760 203024 7812
rect 350632 7760 350684 7812
rect 462780 7760 462832 7812
rect 26516 7692 26568 7744
rect 200304 7692 200356 7744
rect 229836 7692 229888 7744
rect 270592 7692 270644 7744
rect 299572 7692 299624 7744
rect 313832 7692 313884 7744
rect 353392 7692 353444 7744
rect 473452 7692 473504 7744
rect 21824 7624 21876 7676
rect 198832 7624 198884 7676
rect 222752 7624 222804 7676
rect 267924 7624 267976 7676
rect 305000 7624 305052 7676
rect 331588 7624 331640 7676
rect 333244 7624 333296 7676
rect 345756 7624 345808 7676
rect 354772 7624 354824 7676
rect 476948 7624 477000 7676
rect 4068 7556 4120 7608
rect 193312 7556 193364 7608
rect 213368 7556 213420 7608
rect 264244 7556 264296 7608
rect 313280 7556 313332 7608
rect 354036 7556 354088 7608
rect 360200 7556 360252 7608
rect 492312 7556 492364 7608
rect 3424 6808 3476 6860
rect 189724 6808 189776 6860
rect 246396 6400 246448 6452
rect 276112 6400 276164 6452
rect 242992 6332 243044 6384
rect 274916 6332 274968 6384
rect 309140 6332 309192 6384
rect 343364 6332 343416 6384
rect 207388 6264 207440 6316
rect 247684 6264 247736 6316
rect 332600 6264 332652 6316
rect 413100 6264 413152 6316
rect 205088 6196 205140 6248
rect 253204 6196 253256 6248
rect 300952 6196 301004 6248
rect 317328 6196 317380 6248
rect 335360 6196 335412 6248
rect 420184 6196 420236 6248
rect 65524 6128 65576 6180
rect 214104 6128 214156 6180
rect 227536 6128 227588 6180
rect 269304 6128 269356 6180
rect 303620 6128 303672 6180
rect 325608 6128 325660 6180
rect 336740 6128 336792 6180
rect 423772 6128 423824 6180
rect 390560 5176 390612 5228
rect 390928 5176 390980 5228
rect 367100 5108 367152 5160
rect 512460 5108 512512 5160
rect 54944 5040 54996 5092
rect 209872 5040 209924 5092
rect 372712 5040 372764 5092
rect 526628 5040 526680 5092
rect 12348 4972 12400 5024
rect 195980 4972 196032 5024
rect 218152 4972 218204 5024
rect 235264 4972 235316 5024
rect 249984 4972 250036 5024
rect 277676 4972 277728 5024
rect 372620 4972 372672 5024
rect 530124 4972 530176 5024
rect 2872 4904 2924 4956
rect 191840 4904 191892 4956
rect 235816 4904 235868 4956
rect 271972 4904 272024 4956
rect 306380 4904 306432 4956
rect 336280 4904 336332 4956
rect 374000 4904 374052 4956
rect 533712 4904 533764 4956
rect 1676 4836 1728 4888
rect 192024 4836 192076 4888
rect 201500 4836 201552 4888
rect 260840 4836 260892 4888
rect 318800 4836 318852 4888
rect 370596 4836 370648 4888
rect 376760 4836 376812 4888
rect 540796 4836 540848 4888
rect 572 4768 624 4820
rect 191932 4768 191984 4820
rect 195612 4768 195664 4820
rect 257344 4768 257396 4820
rect 320180 4768 320232 4820
rect 374092 4768 374144 4820
rect 378140 4768 378192 4820
rect 544384 4768 544436 4820
rect 300124 4496 300176 4548
rect 306748 4496 306800 4548
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 347044 4156 347096 4208
rect 352840 4156 352892 4208
rect 46664 4088 46716 4140
rect 207020 4088 207072 4140
rect 265348 4088 265400 4140
rect 282920 4088 282972 4140
rect 285404 4088 285456 4140
rect 289084 4088 289136 4140
rect 345020 4088 345072 4140
rect 447416 4088 447468 4140
rect 43076 4020 43128 4072
rect 205640 4020 205692 4072
rect 262956 4020 263008 4072
rect 281632 4020 281684 4072
rect 283104 4020 283156 4072
rect 288532 4020 288584 4072
rect 347780 4020 347832 4072
rect 454500 4020 454552 4072
rect 39580 3952 39632 4004
rect 204536 3952 204588 4004
rect 259552 3952 259604 4004
rect 280344 3952 280396 4004
rect 280712 3952 280764 4004
rect 287244 3952 287296 4004
rect 295984 3952 296036 4004
rect 299664 3952 299716 4004
rect 349252 3952 349304 4004
rect 458088 3952 458140 4004
rect 35992 3884 36044 3936
rect 204352 3884 204404 3936
rect 255872 3884 255924 3936
rect 278872 3884 278924 3936
rect 295340 3884 295392 3936
rect 301964 3884 302016 3936
rect 349160 3884 349212 3936
rect 461584 3884 461636 3936
rect 32404 3816 32456 3868
rect 202880 3816 202932 3868
rect 252376 3816 252428 3868
rect 277584 3816 277636 3868
rect 350540 3816 350592 3868
rect 465172 3816 465224 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 28908 3748 28960 3800
rect 201776 3748 201828 3800
rect 248788 3748 248840 3800
rect 277492 3748 277544 3800
rect 296812 3748 296864 3800
rect 309048 3748 309100 3800
rect 351920 3748 351972 3800
rect 468668 3748 468720 3800
rect 25320 3680 25372 3732
rect 200212 3680 200264 3732
rect 245200 3680 245252 3732
rect 276204 3680 276256 3732
rect 293960 3680 294012 3732
rect 297272 3680 297324 3732
rect 14740 3612 14792 3664
rect 21364 3612 21416 3664
rect 24216 3612 24268 3664
rect 200120 3612 200172 3664
rect 241704 3612 241756 3664
rect 274732 3612 274784 3664
rect 276020 3612 276072 3664
rect 285864 3612 285916 3664
rect 296720 3612 296772 3664
rect 298100 3612 298152 3664
rect 353300 3680 353352 3732
rect 472256 3680 472308 3732
rect 19432 3544 19484 3596
rect 197636 3544 197688 3596
rect 238116 3544 238168 3596
rect 273536 3544 273588 3596
rect 277124 3544 277176 3596
rect 287152 3544 287204 3596
rect 290188 3544 290240 3596
rect 291292 3544 291344 3596
rect 292580 3544 292632 3596
rect 293316 3544 293368 3596
rect 295432 3544 295484 3596
rect 304356 3544 304408 3596
rect 307944 3612 307996 3664
rect 354680 3612 354732 3664
rect 475752 3612 475804 3664
rect 312636 3544 312688 3596
rect 356060 3544 356112 3596
rect 17040 3476 17092 3528
rect 18604 3476 18656 3528
rect 20628 3476 20680 3528
rect 198740 3476 198792 3528
rect 218060 3476 218112 3528
rect 219256 3476 219308 3528
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 259460 3476 259512 3528
rect 260656 3476 260708 3528
rect 272432 3476 272484 3528
rect 284392 3476 284444 3528
rect 294052 3476 294104 3528
rect 298468 3476 298520 3528
rect 299480 3476 299532 3528
rect 316224 3476 316276 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 357532 3476 357584 3528
rect 358728 3476 358780 3528
rect 390744 3544 390796 3596
rect 582196 3544 582248 3596
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 547880 3476 547932 3528
rect 548708 3476 548760 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 570604 3476 570656 3528
rect 571524 3476 571576 3528
rect 571984 3476 572036 3528
rect 572720 3476 572772 3528
rect 6460 3408 6512 3460
rect 10324 3408 10376 3460
rect 15936 3408 15988 3460
rect 17224 3408 17276 3460
rect 11152 3340 11204 3392
rect 194784 3408 194836 3460
rect 231032 3408 231084 3460
rect 270868 3408 270920 3460
rect 273628 3408 273680 3460
rect 285772 3408 285824 3460
rect 300860 3408 300912 3460
rect 319720 3408 319772 3460
rect 365720 3408 365772 3460
rect 367008 3408 367060 3460
rect 390560 3408 390612 3460
rect 581000 3408 581052 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 106924 3340 106976 3392
rect 227720 3340 227772 3392
rect 266544 3340 266596 3392
rect 283012 3340 283064 3392
rect 296904 3340 296956 3392
rect 305552 3340 305604 3392
rect 342260 3340 342312 3392
rect 440240 3340 440292 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 572076 3340 572128 3392
rect 573916 3340 573968 3392
rect 114008 3272 114060 3324
rect 230480 3272 230532 3324
rect 268844 3272 268896 3324
rect 284300 3272 284352 3324
rect 339500 3272 339552 3324
rect 433248 3272 433300 3324
rect 121092 3204 121144 3256
rect 233240 3204 233292 3256
rect 270040 3204 270092 3256
rect 284484 3204 284536 3256
rect 297364 3204 297416 3256
rect 300768 3204 300820 3256
rect 338120 3204 338172 3256
rect 234620 3136 234672 3188
rect 272064 3136 272116 3188
rect 292856 3136 292908 3188
rect 296076 3136 296128 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 407120 3136 407172 3188
rect 408408 3136 408460 3188
rect 415400 3204 415452 3256
rect 416688 3204 416740 3256
rect 423680 3204 423732 3256
rect 424968 3204 425020 3256
rect 426164 3136 426216 3188
rect 284300 3000 284352 3052
rect 288624 3000 288676 3052
rect 292764 3000 292816 3052
rect 294880 3000 294932 3052
rect 9956 2864 10008 2916
rect 14464 2864 14516 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3332 632120 3384 632126
rect 3330 632088 3332 632097
rect 3384 632088 3386 632097
rect 3330 632023 3386 632032
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 605946 2820 606047
rect 2780 605940 2832 605946
rect 2780 605882 2832 605888
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501362 3372 501735
rect 3332 501356 3384 501362
rect 3332 501298 3384 501304
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3436 380866 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3424 380860 3476 380866
rect 3424 380802 3476 380808
rect 3528 373998 3556 658135
rect 4804 605940 4856 605946
rect 4804 605882 4856 605888
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 373992 3568 373998
rect 3516 373934 3568 373940
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 267714 3464 371311
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3424 267708 3476 267714
rect 3424 267650 3476 267656
rect 3528 260846 3556 358391
rect 3620 340882 3648 566879
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3608 340876 3660 340882
rect 3608 340818 3660 340824
rect 3712 333946 3740 553823
rect 3790 462632 3846 462641
rect 3790 462567 3846 462576
rect 3700 333940 3752 333946
rect 3700 333882 3752 333888
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3516 260840 3568 260846
rect 3516 260782 3568 260788
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 220794 3464 254079
rect 3620 247042 3648 319223
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3608 247036 3660 247042
rect 3608 246978 3660 246984
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3424 220788 3476 220794
rect 3424 220730 3476 220736
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 206990 3464 214911
rect 3528 213926 3556 241023
rect 3712 240106 3740 306167
rect 3804 300830 3832 462567
rect 3882 449576 3938 449585
rect 3882 449511 3938 449520
rect 3792 300824 3844 300830
rect 3792 300766 3844 300772
rect 3896 293962 3924 449511
rect 3974 423600 4030 423609
rect 3974 423535 4030 423544
rect 3884 293956 3936 293962
rect 3884 293898 3936 293904
rect 3790 293176 3846 293185
rect 3790 293111 3846 293120
rect 3700 240100 3752 240106
rect 3700 240042 3752 240048
rect 3804 234598 3832 293111
rect 3988 287026 4016 423535
rect 4816 353258 4844 605882
rect 6932 392630 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 18604 683188 18656 683194
rect 18604 683130 18656 683136
rect 13084 618316 13136 618322
rect 13084 618258 13136 618264
rect 8944 501356 8996 501362
rect 8944 501298 8996 501304
rect 6920 392624 6972 392630
rect 6920 392566 6972 392572
rect 4804 353252 4856 353258
rect 4804 353194 4856 353200
rect 4066 345400 4122 345409
rect 4066 345335 4122 345344
rect 3976 287020 4028 287026
rect 3976 286962 4028 286968
rect 3882 267200 3938 267209
rect 3882 267135 3938 267144
rect 3792 234592 3844 234598
rect 3792 234534 3844 234540
rect 3896 227730 3924 267135
rect 4080 253910 4108 345335
rect 8956 314634 8984 501298
rect 10324 397520 10376 397526
rect 10324 397462 10376 397468
rect 8944 314628 8996 314634
rect 8944 314570 8996 314576
rect 10336 274650 10364 397462
rect 13096 360194 13124 618258
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 13084 360188 13136 360194
rect 13084 360130 13136 360136
rect 14476 320142 14504 514762
rect 17224 409896 17276 409902
rect 17224 409838 17276 409844
rect 14464 320136 14516 320142
rect 14464 320078 14516 320084
rect 17236 280158 17264 409838
rect 18616 387802 18644 683130
rect 21364 632120 21416 632126
rect 21364 632062 21416 632068
rect 18604 387796 18656 387802
rect 18604 387738 18656 387744
rect 21376 367062 21404 632062
rect 22744 579692 22796 579698
rect 22744 579634 22796 579640
rect 21364 367056 21416 367062
rect 21364 366998 21416 367004
rect 22756 347750 22784 579634
rect 23492 392698 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 26884 527196 26936 527202
rect 26884 527138 26936 527144
rect 23480 392692 23532 392698
rect 23480 392634 23532 392640
rect 22744 347744 22796 347750
rect 22744 347686 22796 347692
rect 26896 327078 26924 527138
rect 32404 474768 32456 474774
rect 32404 474710 32456 474716
rect 26884 327072 26936 327078
rect 26884 327014 26936 327020
rect 32416 307766 32444 474710
rect 40052 392766 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 392834 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 392902 88380 702406
rect 104912 392970 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 393038 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 393106 153240 702406
rect 169772 393174 169800 702406
rect 169760 393168 169812 393174
rect 169760 393110 169812 393116
rect 153200 393100 153252 393106
rect 153200 393042 153252 393048
rect 136640 393032 136692 393038
rect 136640 392974 136692 392980
rect 104900 392964 104952 392970
rect 104900 392906 104952 392912
rect 88340 392896 88392 392902
rect 88340 392838 88392 392844
rect 71780 392828 71832 392834
rect 71780 392770 71832 392776
rect 40040 392760 40092 392766
rect 40040 392702 40092 392708
rect 201512 392630 201540 702986
rect 217876 392828 217928 392834
rect 217876 392770 217928 392776
rect 210516 392760 210568 392766
rect 210516 392702 210568 392708
rect 203064 392692 203116 392698
rect 203064 392634 203116 392640
rect 195704 392624 195756 392630
rect 195704 392566 195756 392572
rect 201500 392624 201552 392630
rect 201500 392566 201552 392572
rect 195716 389980 195744 392566
rect 203076 389980 203104 392634
rect 210528 389980 210556 392702
rect 217888 389980 217916 392770
rect 218072 392698 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 232688 392964 232740 392970
rect 232688 392906 232740 392912
rect 225328 392896 225380 392902
rect 225328 392838 225380 392844
rect 218060 392692 218112 392698
rect 218060 392634 218112 392640
rect 225340 389980 225368 392838
rect 232700 389980 232728 392906
rect 234632 392766 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 254952 393168 255004 393174
rect 254952 393110 255004 393116
rect 247500 393100 247552 393106
rect 247500 393042 247552 393048
rect 240140 393032 240192 393038
rect 240140 392974 240192 392980
rect 234620 392760 234672 392766
rect 234620 392702 234672 392708
rect 240152 389980 240180 392974
rect 247512 389980 247540 393042
rect 254964 389980 254992 393110
rect 266372 392630 266400 697546
rect 277124 392760 277176 392766
rect 277124 392702 277176 392708
rect 269764 392692 269816 392698
rect 269764 392634 269816 392640
rect 262312 392624 262364 392630
rect 262312 392566 262364 392572
rect 266360 392624 266412 392630
rect 266360 392566 266412 392572
rect 262324 389980 262352 392566
rect 269776 389980 269804 392634
rect 277136 389980 277164 392702
rect 282932 392698 282960 702406
rect 299492 393314 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 328460 700868 328512 700874
rect 328460 700810 328512 700816
rect 306380 700460 306432 700466
rect 306380 700402 306432 700408
rect 299400 393286 299520 393314
rect 282920 392692 282972 392698
rect 282920 392634 282972 392640
rect 291936 392692 291988 392698
rect 291936 392634 291988 392640
rect 284576 392624 284628 392630
rect 284576 392566 284628 392572
rect 284588 389980 284616 392566
rect 291948 389980 291976 392634
rect 299400 389980 299428 393286
rect 306392 389994 306420 700402
rect 313280 700392 313332 700398
rect 313280 700334 313332 700340
rect 313292 402974 313320 700334
rect 321560 700324 321612 700330
rect 321560 700266 321612 700272
rect 313292 402946 313872 402974
rect 313844 389994 313872 402946
rect 306392 389966 306774 389994
rect 313844 389966 314226 389994
rect 321572 389980 321600 700266
rect 328472 402974 328500 700810
rect 332520 700466 332548 703520
rect 335360 700800 335412 700806
rect 335360 700742 335412 700748
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 335372 402974 335400 700742
rect 343640 700732 343692 700738
rect 343640 700674 343692 700680
rect 328472 402946 328592 402974
rect 335372 402946 335952 402974
rect 328564 389994 328592 402946
rect 335924 389994 335952 402946
rect 343652 389994 343680 700674
rect 348804 700398 348832 703520
rect 350540 700664 350592 700670
rect 350540 700606 350592 700612
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 350552 402974 350580 700606
rect 357440 700596 357492 700602
rect 357440 700538 357492 700544
rect 357452 402974 357480 700538
rect 364996 700330 365024 703520
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 413664 700806 413692 703520
rect 413652 700800 413704 700806
rect 413652 700742 413704 700748
rect 429856 700738 429884 703520
rect 429844 700732 429896 700738
rect 429844 700674 429896 700680
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 494808 700534 494836 703520
rect 365720 700528 365772 700534
rect 365720 700470 365772 700476
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 350552 402946 350856 402974
rect 357452 402946 358216 402974
rect 350828 389994 350856 402946
rect 358188 389994 358216 402946
rect 365732 389994 365760 700470
rect 527192 700466 527220 703520
rect 372620 700460 372672 700466
rect 372620 700402 372672 700408
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 372632 402974 372660 700402
rect 543476 700398 543504 703520
rect 379520 700392 379572 700398
rect 379520 700334 379572 700340
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 379532 402974 379560 700334
rect 559668 700330 559696 703520
rect 387800 700324 387852 700330
rect 387800 700266 387852 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 372632 402946 373120 402974
rect 379532 402946 380480 402974
rect 373092 389994 373120 402946
rect 380452 389994 380480 402946
rect 387812 389994 387840 700266
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 406384 683188 406436 683194
rect 406384 683130 406436 683136
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 395344 670744 395396 670750
rect 395344 670686 395396 670692
rect 393964 630692 394016 630698
rect 393964 630634 394016 630640
rect 328564 389966 329038 389994
rect 335924 389966 336398 389994
rect 343652 389966 343850 389994
rect 350828 389966 351210 389994
rect 358188 389966 358662 389994
rect 365732 389966 366022 389994
rect 373092 389966 373474 389994
rect 380452 389966 380834 389994
rect 387812 389966 388286 389994
rect 189080 387796 189132 387802
rect 189080 387738 189132 387744
rect 189092 386617 189120 387738
rect 189078 386608 189134 386617
rect 189078 386543 189134 386552
rect 189080 380860 189132 380866
rect 189080 380802 189132 380808
rect 189092 379953 189120 380802
rect 189078 379944 189134 379953
rect 189078 379879 189134 379888
rect 189080 373992 189132 373998
rect 189080 373934 189132 373940
rect 189092 373289 189120 373934
rect 189078 373280 189134 373289
rect 189078 373215 189134 373224
rect 393872 368144 393924 368150
rect 393870 368112 393872 368121
rect 393924 368112 393926 368121
rect 393870 368047 393926 368056
rect 189080 367056 189132 367062
rect 189080 366998 189132 367004
rect 189092 366625 189120 366998
rect 189078 366616 189134 366625
rect 189078 366551 189134 366560
rect 393976 362001 394004 630634
rect 394516 387796 394568 387802
rect 394516 387738 394568 387744
rect 394528 386889 394556 387738
rect 394514 386880 394570 386889
rect 394514 386815 394570 386824
rect 394608 380860 394660 380866
rect 394608 380802 394660 380808
rect 394620 380633 394648 380802
rect 394606 380624 394662 380633
rect 394606 380559 394662 380568
rect 395356 375358 395384 670686
rect 400864 643136 400916 643142
rect 400864 643078 400916 643084
rect 399484 536852 399536 536858
rect 399484 536794 399536 536800
rect 396724 404388 396776 404394
rect 396724 404330 396776 404336
rect 394148 375352 394200 375358
rect 394148 375294 394200 375300
rect 395344 375352 395396 375358
rect 395344 375294 395396 375300
rect 394160 374377 394188 375294
rect 394146 374368 394202 374377
rect 394146 374303 394202 374312
rect 394056 364404 394108 364410
rect 394056 364346 394108 364352
rect 393962 361992 394018 362001
rect 393962 361927 394018 361936
rect 189080 360188 189132 360194
rect 189080 360130 189132 360136
rect 189092 359961 189120 360130
rect 189078 359952 189134 359961
rect 189078 359887 189134 359896
rect 189078 353288 189134 353297
rect 189078 353223 189080 353232
rect 189132 353223 189134 353232
rect 189080 353194 189132 353200
rect 189080 347744 189132 347750
rect 189080 347686 189132 347692
rect 189092 346633 189120 347686
rect 189078 346624 189134 346633
rect 189078 346559 189134 346568
rect 189080 340876 189132 340882
rect 189080 340818 189132 340824
rect 189092 339969 189120 340818
rect 189078 339960 189134 339969
rect 189078 339895 189134 339904
rect 189080 333940 189132 333946
rect 189080 333882 189132 333888
rect 189092 333305 189120 333882
rect 189078 333296 189134 333305
rect 189078 333231 189134 333240
rect 393964 331220 394016 331226
rect 393964 331162 394016 331168
rect 393976 330857 394004 331162
rect 393962 330848 394018 330857
rect 393962 330783 394018 330792
rect 189080 327072 189132 327078
rect 189080 327014 189132 327020
rect 189092 326641 189120 327014
rect 189078 326632 189134 326641
rect 189078 326567 189134 326576
rect 189080 320136 189132 320142
rect 189080 320078 189132 320084
rect 189092 319977 189120 320078
rect 189078 319968 189134 319977
rect 189078 319903 189134 319912
rect 189080 314628 189132 314634
rect 189080 314570 189132 314576
rect 189092 313313 189120 314570
rect 189078 313304 189134 313313
rect 189078 313239 189134 313248
rect 393964 311908 394016 311914
rect 393964 311850 394016 311856
rect 32404 307760 32456 307766
rect 32404 307702 32456 307708
rect 189080 307760 189132 307766
rect 189080 307702 189132 307708
rect 189092 306649 189120 307702
rect 189078 306640 189134 306649
rect 189078 306575 189134 306584
rect 189080 300824 189132 300830
rect 189080 300766 189132 300772
rect 189092 299985 189120 300766
rect 189078 299976 189134 299985
rect 189078 299911 189134 299920
rect 189080 293956 189132 293962
rect 189080 293898 189132 293904
rect 189092 293321 189120 293898
rect 189078 293312 189134 293321
rect 189078 293247 189134 293256
rect 189080 287020 189132 287026
rect 189080 286962 189132 286968
rect 189092 286657 189120 286962
rect 189078 286648 189134 286657
rect 189078 286583 189134 286592
rect 393688 281308 393740 281314
rect 393688 281250 393740 281256
rect 393700 281081 393728 281250
rect 393686 281072 393742 281081
rect 393686 281007 393742 281016
rect 17224 280152 17276 280158
rect 17224 280094 17276 280100
rect 189080 280152 189132 280158
rect 189080 280094 189132 280100
rect 189092 279993 189120 280094
rect 189078 279984 189134 279993
rect 189078 279919 189134 279928
rect 10324 274644 10376 274650
rect 10324 274586 10376 274592
rect 189080 274644 189132 274650
rect 189080 274586 189132 274592
rect 189092 273329 189120 274586
rect 189078 273320 189134 273329
rect 189078 273255 189134 273264
rect 189080 267708 189132 267714
rect 189080 267650 189132 267656
rect 189092 266665 189120 267650
rect 189078 266656 189134 266665
rect 189078 266591 189134 266600
rect 189080 260840 189132 260846
rect 189080 260782 189132 260788
rect 189092 260001 189120 260782
rect 189078 259992 189134 260001
rect 189078 259927 189134 259936
rect 4068 253904 4120 253910
rect 4068 253846 4120 253852
rect 189080 253904 189132 253910
rect 189080 253846 189132 253852
rect 189092 253337 189120 253846
rect 189078 253328 189134 253337
rect 189078 253263 189134 253272
rect 393976 249937 394004 311850
rect 394068 268569 394096 364346
rect 394608 356040 394660 356046
rect 394608 355982 394660 355988
rect 394620 355745 394648 355982
rect 394606 355736 394662 355745
rect 394606 355671 394662 355680
rect 394608 350532 394660 350538
rect 394608 350474 394660 350480
rect 394620 349489 394648 350474
rect 394606 349480 394662 349489
rect 394606 349415 394662 349424
rect 394240 343596 394292 343602
rect 394240 343538 394292 343544
rect 394252 343233 394280 343538
rect 394238 343224 394294 343233
rect 394238 343159 394294 343168
rect 394608 338088 394660 338094
rect 394608 338030 394660 338036
rect 394620 337113 394648 338030
rect 394606 337104 394662 337113
rect 394606 337039 394662 337048
rect 394608 325644 394660 325650
rect 394608 325586 394660 325592
rect 394620 324601 394648 325586
rect 394606 324592 394662 324601
rect 394606 324527 394662 324536
rect 394608 318776 394660 318782
rect 394608 318718 394660 318724
rect 394620 318345 394648 318718
rect 394606 318336 394662 318345
rect 394606 318271 394662 318280
rect 394608 313268 394660 313274
rect 394608 313210 394660 313216
rect 394620 312225 394648 313210
rect 394606 312216 394662 312225
rect 394606 312151 394662 312160
rect 394240 306332 394292 306338
rect 394240 306274 394292 306280
rect 394252 305969 394280 306274
rect 394238 305960 394294 305969
rect 394238 305895 394294 305904
rect 394608 300824 394660 300830
rect 394608 300766 394660 300772
rect 394620 299713 394648 300766
rect 394606 299704 394662 299713
rect 394606 299639 394662 299648
rect 394608 293956 394660 293962
rect 394608 293898 394660 293904
rect 394620 293457 394648 293898
rect 394606 293448 394662 293457
rect 394606 293383 394662 293392
rect 394608 288380 394660 288386
rect 394608 288322 394660 288328
rect 394620 287337 394648 288322
rect 394606 287328 394662 287337
rect 394606 287263 394662 287272
rect 396736 281314 396764 404330
rect 399496 331226 399524 536794
rect 400876 368150 400904 643078
rect 405004 576904 405056 576910
rect 405004 576846 405056 576852
rect 403624 470620 403676 470626
rect 403624 470562 403676 470568
rect 400864 368144 400916 368150
rect 400864 368086 400916 368092
rect 399484 331220 399536 331226
rect 399484 331162 399536 331168
rect 403636 306338 403664 470562
rect 405016 343602 405044 576846
rect 406396 380866 406424 683130
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 579986 577688 580042 577697
rect 579986 577623 580042 577632
rect 580000 576910 580028 577623
rect 579988 576904 580040 576910
rect 579988 576846 580040 576852
rect 579618 537840 579674 537849
rect 579618 537775 579674 537784
rect 579632 536858 579660 537775
rect 579620 536852 579672 536858
rect 579620 536794 579672 536800
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 549904 456816 549956 456822
rect 549904 456758 549956 456764
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 407764 418192 407816 418198
rect 407764 418134 407816 418140
rect 406384 380860 406436 380866
rect 406384 380802 406436 380808
rect 405004 343596 405056 343602
rect 405004 343538 405056 343544
rect 403624 306332 403676 306338
rect 403624 306274 403676 306280
rect 407776 288386 407804 418134
rect 549916 300830 549944 456758
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580276 387802 580304 697167
rect 580354 617536 580410 617545
rect 580354 617471 580410 617480
rect 580264 387796 580316 387802
rect 580264 387738 580316 387744
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 549904 300824 549956 300830
rect 549904 300766 549956 300772
rect 407764 288380 407816 288386
rect 407764 288322 407816 288328
rect 396724 281308 396776 281314
rect 396724 281250 396776 281256
rect 580276 276010 580304 378383
rect 580368 356046 580396 617471
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580356 356040 580408 356046
rect 580356 355982 580408 355988
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 394608 276004 394660 276010
rect 394608 275946 394660 275952
rect 580264 276004 580316 276010
rect 580264 275946 580316 275952
rect 394620 274825 394648 275946
rect 394606 274816 394662 274825
rect 394606 274751 394662 274760
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 394054 268560 394110 268569
rect 394054 268495 394110 268504
rect 394608 263560 394660 263566
rect 394608 263502 394660 263508
rect 394620 262449 394648 263502
rect 394606 262440 394662 262449
rect 394606 262375 394662 262384
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 394056 258120 394108 258126
rect 394056 258062 394108 258068
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 393962 249928 394018 249937
rect 393962 249863 394018 249872
rect 189080 247036 189132 247042
rect 189080 246978 189132 246984
rect 189092 246673 189120 246978
rect 189078 246664 189134 246673
rect 189078 246599 189134 246608
rect 189080 240100 189132 240106
rect 189080 240042 189132 240048
rect 189092 240009 189120 240042
rect 189078 240000 189134 240009
rect 189078 239935 189134 239944
rect 189080 234592 189132 234598
rect 189080 234534 189132 234540
rect 189092 233345 189120 234534
rect 189078 233336 189134 233345
rect 189078 233271 189134 233280
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 3884 227724 3936 227730
rect 3884 227666 3936 227672
rect 189080 227724 189132 227730
rect 189080 227666 189132 227672
rect 189092 226681 189120 227666
rect 189078 226672 189134 226681
rect 189078 226607 189134 226616
rect 189080 220788 189132 220794
rect 189080 220730 189132 220736
rect 189092 220017 189120 220730
rect 189078 220008 189134 220017
rect 189078 219943 189134 219952
rect 393976 218793 394004 231814
rect 394068 231305 394096 258062
rect 394608 256692 394660 256698
rect 394608 256634 394660 256640
rect 394620 256193 394648 256634
rect 394606 256184 394662 256193
rect 394606 256119 394662 256128
rect 394608 244248 394660 244254
rect 394608 244190 394660 244196
rect 394620 243681 394648 244190
rect 394606 243672 394662 243681
rect 394606 243607 394662 243616
rect 580276 238746 580304 272167
rect 580368 263566 580396 351863
rect 580460 350538 580488 590951
rect 580538 564360 580594 564369
rect 580538 564295 580594 564304
rect 580448 350532 580500 350538
rect 580448 350474 580500 350480
rect 580552 338094 580580 564295
rect 580630 524512 580686 524521
rect 580630 524447 580686 524456
rect 580540 338088 580592 338094
rect 580540 338030 580592 338036
rect 580644 325650 580672 524447
rect 580722 511320 580778 511329
rect 580722 511255 580778 511264
rect 580632 325644 580684 325650
rect 580632 325586 580684 325592
rect 580446 325272 580502 325281
rect 580446 325207 580502 325216
rect 580356 263560 580408 263566
rect 580356 263502 580408 263508
rect 580460 256698 580488 325207
rect 580736 318782 580764 511255
rect 580814 484664 580870 484673
rect 580814 484599 580870 484608
rect 580724 318776 580776 318782
rect 580724 318718 580776 318724
rect 580828 313274 580856 484599
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580816 313268 580868 313274
rect 580816 313210 580868 313216
rect 580538 298752 580594 298761
rect 580538 298687 580594 298696
rect 580448 256692 580500 256698
rect 580448 256634 580500 256640
rect 580354 245576 580410 245585
rect 580354 245511 580410 245520
rect 394608 238740 394660 238746
rect 394608 238682 394660 238688
rect 580264 238740 580316 238746
rect 580264 238682 580316 238688
rect 394620 237561 394648 238682
rect 394606 237552 394662 237561
rect 394606 237487 394662 237496
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 394054 231296 394110 231305
rect 394054 231231 394110 231240
rect 580368 226302 580396 245511
rect 580552 244254 580580 298687
rect 580920 293962 580948 431559
rect 580908 293956 580960 293962
rect 580908 293898 580960 293904
rect 580540 244248 580592 244254
rect 580540 244190 580592 244196
rect 394608 226296 394660 226302
rect 394608 226238 394660 226244
rect 580356 226296 580408 226302
rect 580356 226238 580408 226244
rect 394620 225049 394648 226238
rect 394606 225040 394662 225049
rect 394606 224975 394662 224984
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 393962 218784 394018 218793
rect 393962 218719 394018 218728
rect 580184 218074 580212 218991
rect 393964 218068 394016 218074
rect 393964 218010 394016 218016
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 3516 213920 3568 213926
rect 3516 213862 3568 213868
rect 189080 213920 189132 213926
rect 189080 213862 189132 213868
rect 189092 213353 189120 213862
rect 189078 213344 189134 213353
rect 189078 213279 189134 213288
rect 393976 212673 394004 218010
rect 393962 212664 394018 212673
rect 393962 212599 394018 212608
rect 3424 206984 3476 206990
rect 3424 206926 3476 206932
rect 189080 206984 189132 206990
rect 189080 206926 189132 206932
rect 189092 206689 189120 206926
rect 189078 206680 189134 206689
rect 189078 206615 189134 206624
rect 394606 206408 394662 206417
rect 394606 206343 394662 206352
rect 394620 206310 394648 206343
rect 394608 206304 394660 206310
rect 394608 206246 394660 206252
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 3146 201920 3202 201929
rect 3146 201855 3202 201864
rect 3160 200122 3188 201855
rect 394054 200152 394110 200161
rect 3148 200116 3200 200122
rect 3148 200058 3200 200064
rect 189080 200116 189132 200122
rect 394054 200087 394110 200096
rect 189080 200058 189132 200064
rect 189092 200025 189120 200058
rect 189078 200016 189134 200025
rect 189078 199951 189134 199960
rect 393962 193896 394018 193905
rect 393962 193831 394018 193840
rect 189078 193352 189134 193361
rect 189078 193287 189134 193296
rect 189092 193254 189120 193287
rect 3424 193248 3476 193254
rect 3424 193190 3476 193196
rect 189080 193248 189132 193254
rect 189080 193190 189132 193196
rect 3436 188873 3464 193190
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 189814 186688 189870 186697
rect 189814 186623 189870 186632
rect 189078 180024 189134 180033
rect 189078 179959 189134 179968
rect 189092 179450 189120 179959
rect 3424 179444 3476 179450
rect 3424 179386 3476 179392
rect 189080 179444 189132 179450
rect 189080 179386 189132 179392
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 149841 3464 179386
rect 189722 173360 189778 173369
rect 189722 173295 189778 173304
rect 189078 160032 189134 160041
rect 189078 159967 189134 159976
rect 189092 158778 189120 159967
rect 3608 158772 3660 158778
rect 3608 158714 3660 158720
rect 189080 158772 189132 158778
rect 189080 158714 189132 158720
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3516 139460 3568 139466
rect 3516 139402 3568 139408
rect 3424 137964 3476 137970
rect 3424 137906 3476 137912
rect 3436 136785 3464 137906
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3424 118720 3476 118726
rect 3424 118662 3476 118668
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 118662
rect 3528 58585 3556 139402
rect 3620 97617 3648 158714
rect 189078 140040 189134 140049
rect 189078 139975 189134 139984
rect 189092 139466 189120 139975
rect 189080 139460 189132 139466
rect 189080 139402 189132 139408
rect 189736 137970 189764 173295
rect 189828 164218 189856 186623
rect 393976 179382 394004 193831
rect 394068 193186 394096 200087
rect 394056 193180 394108 193186
rect 394056 193122 394108 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 394238 187776 394294 187785
rect 394238 187711 394294 187720
rect 394146 181520 394202 181529
rect 394146 181455 394202 181464
rect 393964 179376 394016 179382
rect 393964 179318 394016 179324
rect 394054 175264 394110 175273
rect 394054 175199 394110 175208
rect 393962 169008 394018 169017
rect 393962 168943 394018 168952
rect 190182 166696 190238 166705
rect 190182 166631 190238 166640
rect 189816 164212 189868 164218
rect 189816 164154 189868 164160
rect 190090 153368 190146 153377
rect 190090 153303 190146 153312
rect 189998 146704 190054 146713
rect 189998 146639 190054 146648
rect 189724 137964 189776 137970
rect 189724 137906 189776 137912
rect 189906 133376 189962 133385
rect 189906 133311 189962 133320
rect 189814 126712 189870 126721
rect 189814 126647 189870 126656
rect 189078 120048 189134 120057
rect 189078 119983 189134 119992
rect 189092 118726 189120 119983
rect 189080 118720 189132 118726
rect 189080 118662 189132 118668
rect 189722 113384 189778 113393
rect 189722 113319 189778 113328
rect 188344 108656 188396 108662
rect 188344 108598 188396 108604
rect 124220 108588 124272 108594
rect 124220 108530 124272 108536
rect 117320 108520 117372 108526
rect 117320 108462 117372 108468
rect 110420 108452 110472 108458
rect 110420 108394 110472 108400
rect 17224 108384 17276 108390
rect 17224 108326 17276 108332
rect 10324 108316 10376 108322
rect 10324 108258 10376 108264
rect 6920 98660 6972 98666
rect 6920 98602 6972 98608
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 6932 16574 6960 98602
rect 8300 97300 8352 97306
rect 8300 97242 8352 97248
rect 8312 16574 8340 97242
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 10336 3466 10364 108258
rect 14464 101448 14516 101454
rect 14464 101390 14516 101396
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 480 9996 2858
rect 11164 480 11192 3334
rect 12360 480 12388 4966
rect 13556 480 13584 8910
rect 14476 2922 14504 101390
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14752 480 14780 3606
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 480 15976 3402
rect 17052 480 17080 3470
rect 17236 3466 17264 108326
rect 74540 106956 74592 106962
rect 74540 106898 74592 106904
rect 60740 105596 60792 105602
rect 60740 105538 60792 105544
rect 57980 104168 58032 104174
rect 57980 104110 58032 104116
rect 46940 102808 46992 102814
rect 46940 102750 46992 102756
rect 29000 100020 29052 100026
rect 29000 99962 29052 99968
rect 18604 79348 18656 79354
rect 18604 79290 18656 79296
rect 17960 33788 18012 33794
rect 17960 33730 18012 33736
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 33730
rect 18616 3534 18644 79290
rect 27620 68332 27672 68338
rect 27620 68274 27672 68280
rect 21364 62824 21416 62830
rect 21364 62766 21416 62772
rect 21376 3670 21404 62766
rect 27632 16574 27660 68274
rect 29012 16574 29040 99962
rect 34520 95940 34572 95946
rect 34520 95882 34572 95888
rect 30380 43444 30432 43450
rect 30380 43386 30432 43392
rect 30392 16574 30420 43386
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 22560 13116 22612 13122
rect 22560 13058 22612 13064
rect 21824 7676 21876 7682
rect 21824 7618 21876 7624
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 19444 480 19472 3538
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 480 20668 3470
rect 21836 480 21864 7618
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 13058
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 480 24256 3606
rect 25332 480 25360 3674
rect 26528 480 26556 7686
rect 27724 480 27752 16546
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 33600 7812 33652 7818
rect 33600 7754 33652 7760
rect 32404 3868 32456 3874
rect 32404 3810 32456 3816
rect 32416 480 32444 3810
rect 33612 480 33640 7754
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 95882
rect 35900 91792 35952 91798
rect 35900 91734 35952 91740
rect 35912 16574 35940 91734
rect 44180 72480 44232 72486
rect 44180 72422 44232 72428
rect 41420 69692 41472 69698
rect 41420 69634 41472 69640
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37292 16574 37320 17206
rect 41432 16574 41460 69634
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 41432 16546 41920 16574
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 480 36032 3878
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 40684 9036 40736 9042
rect 40684 8978 40736 8984
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39592 480 39620 3946
rect 40696 480 40724 8978
rect 41892 480 41920 16546
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 44192 3398 44220 72422
rect 46952 16574 46980 102750
rect 48320 90364 48372 90370
rect 48320 90306 48372 90312
rect 48332 16574 48360 90306
rect 56600 82136 56652 82142
rect 56600 82078 56652 82084
rect 52460 75200 52512 75206
rect 52460 75142 52512 75148
rect 49700 73840 49752 73846
rect 49700 73782 49752 73788
rect 49712 16574 49740 73782
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44272 10328 44324 10334
rect 44272 10270 44324 10276
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 10270
rect 46664 4140 46716 4146
rect 46664 4082 46716 4088
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 4082
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51080 15904 51132 15910
rect 51080 15846 51132 15852
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 15846
rect 52472 3398 52500 75142
rect 55220 21412 55272 21418
rect 55220 21354 55272 21360
rect 55232 16574 55260 21354
rect 56612 16574 56640 82078
rect 57992 16574 58020 104110
rect 59360 49020 59412 49026
rect 59360 48962 59412 48968
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52552 10396 52604 10402
rect 52552 10338 52604 10344
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 10338
rect 54944 5092 54996 5098
rect 54944 5034 54996 5040
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 5034
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 48962
rect 60752 3398 60780 105538
rect 62120 89004 62172 89010
rect 62120 88946 62172 88952
rect 60832 29640 60884 29646
rect 60832 29582 60884 29588
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 29582
rect 62132 16574 62160 88946
rect 66260 80708 66312 80714
rect 66260 80650 66312 80656
rect 63500 76560 63552 76566
rect 63500 76502 63552 76508
rect 63512 16574 63540 76502
rect 66272 16574 66300 80650
rect 69020 61396 69072 61402
rect 69020 61338 69072 61344
rect 67640 28280 67692 28286
rect 67640 28222 67692 28228
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 6180 65576 6186
rect 65524 6122 65576 6128
rect 65536 480 65564 6122
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 28222
rect 69032 6914 69060 61338
rect 71780 60036 71832 60042
rect 71780 59978 71832 59984
rect 70400 42084 70452 42090
rect 70400 42026 70452 42032
rect 69112 18624 69164 18630
rect 69112 18566 69164 18572
rect 69124 16574 69152 18566
rect 70412 16574 70440 42026
rect 71792 16574 71820 59978
rect 73160 31068 73212 31074
rect 73160 31010 73212 31016
rect 73172 16574 73200 31010
rect 74552 16574 74580 106898
rect 81440 98728 81492 98734
rect 81440 98670 81492 98676
rect 78680 94512 78732 94518
rect 78680 94454 78732 94460
rect 77300 87644 77352 87650
rect 77300 87586 77352 87592
rect 75920 77988 75972 77994
rect 75920 77930 75972 77936
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 77930
rect 77312 6914 77340 87586
rect 77392 26920 77444 26926
rect 77392 26862 77444 26868
rect 77404 16574 77432 26862
rect 78692 16574 78720 94454
rect 81452 16574 81480 98670
rect 89720 93152 89772 93158
rect 89720 93094 89772 93100
rect 85580 58676 85632 58682
rect 85580 58618 85632 58624
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80888 11756 80940 11762
rect 80888 11698 80940 11704
rect 80900 480 80928 11698
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 84200 11824 84252 11830
rect 84200 11766 84252 11772
rect 83280 7880 83332 7886
rect 83280 7822 83332 7828
rect 83292 480 83320 7822
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 11766
rect 85592 3398 85620 58618
rect 88340 54528 88392 54534
rect 88340 54470 88392 54476
rect 86960 47592 87012 47598
rect 86960 47534 87012 47540
rect 85672 25560 85724 25566
rect 85672 25502 85724 25508
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 25502
rect 86972 16574 87000 47534
rect 88352 16574 88380 54470
rect 89732 16574 89760 93094
rect 92480 84856 92532 84862
rect 92480 84798 92532 84804
rect 91100 66904 91152 66910
rect 91100 66846 91152 66852
rect 91112 16574 91140 66846
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 84798
rect 102140 83496 102192 83502
rect 102140 83438 102192 83444
rect 95240 65544 95292 65550
rect 95240 65486 95292 65492
rect 95252 16574 95280 65486
rect 99380 64184 99432 64190
rect 99380 64126 99432 64132
rect 99392 16574 99420 64126
rect 100760 57248 100812 57254
rect 100760 57190 100812 57196
rect 95252 16546 95832 16574
rect 99392 16546 99880 16574
rect 93860 11892 93912 11898
rect 93860 11834 93912 11840
rect 93872 3398 93900 11834
rect 93952 10464 94004 10470
rect 93952 10406 94004 10412
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 10406
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 98184 11960 98236 11966
rect 98184 11902 98236 11908
rect 97448 10532 97500 10538
rect 97448 10474 97500 10480
rect 97460 480 97488 10474
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 11902
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 57190
rect 102152 6914 102180 83438
rect 102232 53100 102284 53106
rect 102232 53042 102284 53048
rect 102244 16574 102272 53042
rect 102244 16546 103376 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 109040 12096 109092 12102
rect 109040 12038 109092 12044
rect 105728 12028 105780 12034
rect 105728 11970 105780 11976
rect 104072 10600 104124 10606
rect 104072 10542 104124 10548
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 10542
rect 105740 480 105768 11970
rect 108120 10668 108172 10674
rect 108120 10610 108172 10616
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 106936 480 106964 3334
rect 108132 480 108160 10610
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 12038
rect 110432 6914 110460 108394
rect 114560 86284 114612 86290
rect 114560 86226 114612 86232
rect 110512 55888 110564 55894
rect 110512 55830 110564 55836
rect 110524 16574 110552 55830
rect 114572 16574 114600 86226
rect 110524 16546 111656 16574
rect 114572 16546 114784 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 112352 13184 112404 13190
rect 112352 13126 112404 13132
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 13126
rect 114008 3324 114060 3330
rect 114008 3266 114060 3272
rect 114020 480 114048 3266
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116400 13252 116452 13258
rect 116400 13194 116452 13200
rect 116412 480 116440 13194
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 108462
rect 121460 51740 121512 51746
rect 121460 51682 121512 51688
rect 118700 35216 118752 35222
rect 118700 35158 118752 35164
rect 118712 16574 118740 35158
rect 121472 16574 121500 51682
rect 124232 16574 124260 108530
rect 157340 107092 157392 107098
rect 157340 107034 157392 107040
rect 125600 107024 125652 107030
rect 125600 106966 125652 106972
rect 118712 16546 118832 16574
rect 121472 16546 122328 16574
rect 124232 16546 124720 16574
rect 118804 480 118832 16546
rect 119896 13320 119948 13326
rect 119896 13262 119948 13268
rect 119908 480 119936 13262
rect 121092 3256 121144 3262
rect 121092 3198 121144 3204
rect 121104 480 121132 3198
rect 122300 480 122328 16546
rect 123024 13388 123076 13394
rect 123024 13330 123076 13336
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 13330
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 106966
rect 131120 101516 131172 101522
rect 131120 101458 131172 101464
rect 129740 96008 129792 96014
rect 129740 95950 129792 95956
rect 128360 94580 128412 94586
rect 128360 94522 128412 94528
rect 126980 82204 127032 82210
rect 126980 82146 127032 82152
rect 126992 480 127020 82146
rect 127072 39364 127124 39370
rect 127072 39306 127124 39312
rect 127084 16574 127112 39306
rect 128372 16574 128400 94522
rect 129752 16574 129780 95950
rect 131132 16574 131160 101458
rect 151820 100088 151872 100094
rect 151820 100030 151872 100036
rect 142160 97368 142212 97374
rect 142160 97310 142212 97316
rect 132500 93220 132552 93226
rect 132500 93162 132552 93168
rect 132512 16574 132540 93162
rect 135260 91860 135312 91866
rect 135260 91802 135312 91808
rect 133880 76628 133932 76634
rect 133880 76570 133932 76576
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 76570
rect 135272 4214 135300 91802
rect 139400 90432 139452 90438
rect 139400 90374 139452 90380
rect 135352 65612 135404 65618
rect 135352 65554 135404 65560
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 135364 3482 135392 65554
rect 138020 64252 138072 64258
rect 138020 64194 138072 64200
rect 136640 37936 136692 37942
rect 136640 37878 136692 37884
rect 136652 16574 136680 37878
rect 138032 16574 138060 64194
rect 139412 16574 139440 90374
rect 140780 36576 140832 36582
rect 140780 36518 140832 36524
rect 140792 16574 140820 36518
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4150
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 97310
rect 143540 89072 143592 89078
rect 143540 89014 143592 89020
rect 143552 480 143580 89014
rect 146300 87712 146352 87718
rect 146300 87654 146352 87660
rect 144920 50380 144972 50386
rect 144920 50322 144972 50328
rect 143632 46232 143684 46238
rect 143632 46174 143684 46180
rect 143644 16574 143672 46174
rect 144932 16574 144960 50322
rect 146312 16574 146340 87654
rect 150440 86352 150492 86358
rect 150440 86294 150492 86300
rect 147680 75268 147732 75274
rect 147680 75210 147732 75216
rect 147692 16574 147720 75210
rect 149060 53168 149112 53174
rect 149060 53110 149112 53116
rect 149072 16574 149100 53110
rect 150452 16574 150480 86294
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 100030
rect 153200 83564 153252 83570
rect 153200 83506 153252 83512
rect 151912 73908 151964 73914
rect 151912 73850 151964 73856
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 73850
rect 153212 16574 153240 83506
rect 154580 72548 154632 72554
rect 154580 72490 154632 72496
rect 154592 16574 154620 72490
rect 155960 62892 156012 62898
rect 155960 62834 156012 62840
rect 155972 16574 156000 62834
rect 157352 16574 157380 107034
rect 169760 105732 169812 105738
rect 169760 105674 169812 105680
rect 160100 105664 160152 105670
rect 160100 105606 160152 105612
rect 158720 40724 158772 40730
rect 158720 40666 158772 40672
rect 158732 16574 158760 40666
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11694 160140 105606
rect 164240 104236 164292 104242
rect 164240 104178 164292 104184
rect 161480 80776 161532 80782
rect 161480 80718 161532 80724
rect 160192 54596 160244 54602
rect 160192 54538 160244 54544
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 160204 6914 160232 54538
rect 161492 16574 161520 80718
rect 162860 69760 162912 69766
rect 162860 69702 162912 69708
rect 162872 16574 162900 69702
rect 164252 16574 164280 104178
rect 165620 79416 165672 79422
rect 165620 79358 165672 79364
rect 165632 16574 165660 79358
rect 167000 68400 167052 68406
rect 167000 68342 167052 68348
rect 167012 16574 167040 68342
rect 168380 22772 168432 22778
rect 168380 22714 168432 22720
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11630
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 11694 168420 22714
rect 169772 16574 169800 105674
rect 173900 104304 173952 104310
rect 173900 104246 173952 104252
rect 171140 102876 171192 102882
rect 171140 102818 171192 102824
rect 171152 16574 171180 102818
rect 172520 24132 172572 24138
rect 172520 24074 172572 24080
rect 172532 16574 172560 24074
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 168472 14476 168524 14482
rect 168472 14418 168524 14424
rect 168380 11688 168432 11694
rect 168380 11630 168432 11636
rect 168484 6914 168512 14418
rect 169576 11688 169628 11694
rect 169576 11630 169628 11636
rect 168392 6886 168512 6914
rect 168392 480 168420 6886
rect 169588 480 169616 11630
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 104246
rect 187700 102944 187752 102950
rect 187700 102886 187752 102892
rect 175280 101584 175332 101590
rect 175280 101526 175332 101532
rect 175292 16574 175320 101526
rect 178040 100156 178092 100162
rect 178040 100098 178092 100104
rect 176660 42152 176712 42158
rect 176660 42094 176712 42100
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 11694 176700 42094
rect 176752 25628 176804 25634
rect 176752 25570 176804 25576
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 25570
rect 178052 16574 178080 100098
rect 182180 98796 182232 98802
rect 182180 98738 182232 98744
rect 179420 84924 179472 84930
rect 179420 84866 179472 84872
rect 179432 16574 179460 84866
rect 180800 66972 180852 66978
rect 180800 66914 180852 66920
rect 180812 16574 180840 66914
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 98738
rect 184940 97436 184992 97442
rect 184940 97378 184992 97384
rect 183560 78056 183612 78062
rect 183560 77998 183612 78004
rect 183572 16574 183600 77998
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11694 184980 97378
rect 185032 71052 185084 71058
rect 185032 70994 185084 71000
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 70994
rect 186320 26988 186372 26994
rect 186320 26930 186372 26936
rect 186332 16574 186360 26930
rect 186332 16546 186912 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 187712 6914 187740 102886
rect 188356 15910 188384 108598
rect 189080 32428 189132 32434
rect 189080 32370 189132 32376
rect 189092 16574 189120 32370
rect 189092 16546 189304 16574
rect 188344 15904 188396 15910
rect 188344 15846 188396 15852
rect 187712 6886 188568 6914
rect 188540 480 188568 6886
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189736 6866 189764 113319
rect 189828 33114 189856 126647
rect 189920 45558 189948 133311
rect 190012 71738 190040 146639
rect 190104 85542 190132 153303
rect 190196 111790 190224 166631
rect 393778 131744 393834 131753
rect 393778 131679 393834 131688
rect 393792 131170 393820 131679
rect 393780 131164 393832 131170
rect 393780 131106 393832 131112
rect 393976 126954 394004 168943
rect 394068 139398 394096 175199
rect 394160 153202 394188 181455
rect 394252 167006 394280 187711
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 394240 167000 394292 167006
rect 394240 166942 394292 166948
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 394514 162888 394570 162897
rect 394514 162823 394570 162832
rect 394422 156632 394478 156641
rect 394422 156567 394478 156576
rect 394148 153196 394200 153202
rect 394148 153138 394200 153144
rect 394330 150376 394386 150385
rect 394330 150311 394386 150320
rect 394238 144120 394294 144129
rect 394238 144055 394294 144064
rect 394056 139392 394108 139398
rect 394056 139334 394108 139340
rect 394146 138000 394202 138009
rect 394146 137935 394202 137944
rect 393964 126948 394016 126954
rect 393964 126890 394016 126896
rect 394054 125488 394110 125497
rect 394054 125423 394110 125432
rect 393962 119232 394018 119241
rect 393962 119167 394018 119176
rect 190184 111784 190236 111790
rect 190184 111726 190236 111732
rect 215496 110214 215694 110242
rect 225156 110226 225446 110242
rect 224960 110220 225012 110226
rect 191944 110078 192234 110106
rect 192312 110078 192602 110106
rect 192680 110078 192970 110106
rect 193324 110078 193430 110106
rect 193600 110078 193798 110106
rect 191840 106820 191892 106826
rect 191840 106762 191892 106768
rect 190092 85536 190144 85542
rect 190092 85478 190144 85484
rect 190000 71732 190052 71738
rect 190000 71674 190052 71680
rect 189908 45552 189960 45558
rect 189908 45494 189960 45500
rect 189816 33108 189868 33114
rect 189816 33050 189868 33056
rect 190460 28348 190512 28354
rect 190460 28290 190512 28296
rect 189724 6860 189776 6866
rect 189724 6802 189776 6808
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 28290
rect 191852 4962 191880 106762
rect 191840 4956 191892 4962
rect 191840 4898 191892 4904
rect 191944 4826 191972 110078
rect 192312 103514 192340 110078
rect 192680 106826 192708 110078
rect 192668 106820 192720 106826
rect 192668 106762 192720 106768
rect 192036 103486 192340 103514
rect 192036 4894 192064 103486
rect 192116 19984 192168 19990
rect 192116 19926 192168 19932
rect 192024 4888 192076 4894
rect 192024 4830 192076 4836
rect 191932 4820 191984 4826
rect 191932 4762 191984 4768
rect 192128 3482 192156 19926
rect 193324 7614 193352 110078
rect 193404 96076 193456 96082
rect 193404 96018 193456 96024
rect 193312 7608 193364 7614
rect 193312 7550 193364 7556
rect 193416 6914 193444 96018
rect 193496 29708 193548 29714
rect 193496 29650 193548 29656
rect 192036 3454 192156 3482
rect 193232 6886 193444 6914
rect 192036 480 192064 3454
rect 193232 480 193260 6886
rect 193508 3482 193536 29650
rect 193600 3641 193628 110078
rect 194244 108322 194272 110092
rect 194232 108316 194284 108322
rect 194232 108258 194284 108264
rect 193864 107772 193916 107778
rect 193864 107714 193916 107720
rect 193876 97306 193904 107714
rect 194612 107710 194640 110092
rect 194980 107778 195008 110092
rect 195072 110078 195454 110106
rect 195532 110078 195822 110106
rect 195992 110078 196282 110106
rect 196360 110078 196650 110106
rect 196728 110078 197018 110106
rect 194968 107772 195020 107778
rect 194968 107714 195020 107720
rect 193956 107704 194008 107710
rect 193956 107646 194008 107652
rect 194600 107704 194652 107710
rect 194600 107646 194652 107652
rect 193968 98666 193996 107646
rect 195072 106842 195100 110078
rect 194704 106814 195100 106842
rect 194704 101454 194732 106814
rect 195532 103514 195560 110078
rect 194796 103486 195560 103514
rect 194692 101448 194744 101454
rect 194692 101390 194744 101396
rect 193956 98660 194008 98666
rect 193956 98602 194008 98608
rect 193864 97300 193916 97306
rect 193864 97242 193916 97248
rect 193586 3632 193642 3641
rect 193586 3567 193642 3576
rect 193508 3454 194456 3482
rect 194796 3466 194824 103486
rect 195992 5030 196020 110078
rect 196360 106842 196388 110078
rect 196084 106814 196388 106842
rect 196084 8974 196112 106814
rect 196728 103514 196756 110078
rect 197464 108390 197492 110092
rect 197556 110078 197846 110106
rect 198016 110078 198306 110106
rect 198384 110078 198674 110106
rect 198752 110078 199042 110106
rect 199120 110078 199502 110106
rect 199580 110078 199870 110106
rect 200132 110078 200330 110106
rect 200408 110078 200698 110106
rect 200776 110078 201158 110106
rect 201526 110078 201724 110106
rect 197452 108384 197504 108390
rect 197452 108326 197504 108332
rect 197452 106140 197504 106146
rect 197452 106082 197504 106088
rect 196176 103486 196756 103514
rect 196176 62830 196204 103486
rect 196164 62824 196216 62830
rect 196164 62766 196216 62772
rect 197464 33794 197492 106082
rect 197556 79354 197584 110078
rect 198016 106146 198044 110078
rect 198004 106140 198056 106146
rect 198004 106082 198056 106088
rect 198384 103514 198412 110078
rect 197648 103486 198412 103514
rect 197544 79348 197596 79354
rect 197544 79290 197596 79296
rect 197452 33788 197504 33794
rect 197452 33730 197504 33736
rect 197544 33788 197596 33794
rect 197544 33730 197596 33736
rect 196808 15904 196860 15910
rect 196808 15846 196860 15852
rect 196072 8968 196124 8974
rect 196072 8910 196124 8916
rect 195980 5024 196032 5030
rect 195980 4966 196032 4972
rect 195612 4820 195664 4826
rect 195612 4762 195664 4768
rect 194428 480 194456 3454
rect 194784 3460 194836 3466
rect 194784 3402 194836 3408
rect 195624 480 195652 4762
rect 196820 480 196848 15846
rect 197556 3482 197584 33730
rect 197648 3602 197676 103486
rect 197636 3596 197688 3602
rect 197636 3538 197688 3544
rect 198752 3534 198780 110078
rect 199120 106842 199148 110078
rect 198844 106814 199148 106842
rect 198844 7682 198872 106814
rect 199580 103514 199608 110078
rect 198936 103486 199608 103514
rect 198936 13122 198964 103486
rect 199016 43512 199068 43518
rect 199016 43454 199068 43460
rect 199028 16574 199056 43454
rect 199028 16546 199148 16574
rect 198924 13116 198976 13122
rect 198924 13058 198976 13064
rect 198832 7676 198884 7682
rect 198832 7618 198884 7624
rect 198740 3528 198792 3534
rect 197556 3454 197952 3482
rect 198740 3470 198792 3476
rect 197924 480 197952 3454
rect 199120 480 199148 16546
rect 200132 3670 200160 110078
rect 200408 103714 200436 110078
rect 200224 103686 200436 103714
rect 200224 3738 200252 103686
rect 200776 103514 200804 110078
rect 201500 106888 201552 106894
rect 201500 106830 201552 106836
rect 200316 103486 200804 103514
rect 200316 7750 200344 103486
rect 201512 100026 201540 106830
rect 201592 106820 201644 106826
rect 201592 106762 201644 106768
rect 201500 100020 201552 100026
rect 201500 99962 201552 99968
rect 201604 43450 201632 106762
rect 201696 68338 201724 110078
rect 201788 110078 201894 110106
rect 202064 110078 202354 110106
rect 202432 110078 202722 110106
rect 202892 110078 203182 110106
rect 203260 110078 203550 110106
rect 203628 110078 203918 110106
rect 201684 68332 201736 68338
rect 201684 68274 201736 68280
rect 201592 43444 201644 43450
rect 201592 43386 201644 43392
rect 200396 17332 200448 17338
rect 200396 17274 200448 17280
rect 200304 7744 200356 7750
rect 200304 7686 200356 7692
rect 200408 6914 200436 17274
rect 200316 6886 200436 6914
rect 200212 3732 200264 3738
rect 200212 3674 200264 3680
rect 200120 3664 200172 3670
rect 200120 3606 200172 3612
rect 200316 480 200344 6886
rect 201500 4888 201552 4894
rect 201500 4830 201552 4836
rect 201512 480 201540 4830
rect 201788 3806 201816 110078
rect 202064 106894 202092 110078
rect 202052 106888 202104 106894
rect 202052 106830 202104 106836
rect 202432 106826 202460 110078
rect 202420 106820 202472 106826
rect 202420 106762 202472 106768
rect 202696 8968 202748 8974
rect 202696 8910 202748 8916
rect 201776 3800 201828 3806
rect 201776 3742 201828 3748
rect 202708 480 202736 8910
rect 202892 3874 202920 110078
rect 203260 106808 203288 110078
rect 203628 107930 203656 110078
rect 202984 106780 203288 106808
rect 203352 107902 203656 107930
rect 202984 7818 203012 106780
rect 203352 103514 203380 107902
rect 203524 107772 203576 107778
rect 203524 107714 203576 107720
rect 203076 103486 203380 103514
rect 203076 95946 203104 103486
rect 203064 95940 203116 95946
rect 203064 95882 203116 95888
rect 203064 18692 203116 18698
rect 203064 18634 203116 18640
rect 203076 16574 203104 18634
rect 203536 17270 203564 107714
rect 203708 107704 203760 107710
rect 203708 107646 203760 107652
rect 203720 103514 203748 107646
rect 203628 103486 203748 103514
rect 203628 91798 203656 103486
rect 203616 91792 203668 91798
rect 203616 91734 203668 91740
rect 203524 17264 203576 17270
rect 203524 17206 203576 17212
rect 203076 16546 203472 16574
rect 202972 7812 203024 7818
rect 202972 7754 203024 7760
rect 202880 3868 202932 3874
rect 202880 3810 202932 3816
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 204364 3942 204392 110092
rect 204732 107710 204760 110092
rect 205192 107778 205220 110092
rect 205284 110078 205574 110106
rect 205744 110078 205942 110106
rect 206020 110078 206402 110106
rect 206480 110078 206770 110106
rect 207124 110078 207230 110106
rect 207308 110078 207598 110106
rect 207676 110078 207966 110106
rect 205180 107772 205232 107778
rect 205180 107714 205232 107720
rect 204720 107704 204772 107710
rect 204720 107646 204772 107652
rect 205284 103514 205312 110078
rect 205640 104100 205692 104106
rect 205640 104042 205692 104048
rect 204548 103486 205312 103514
rect 204548 4010 204576 103486
rect 205088 6248 205140 6254
rect 205088 6190 205140 6196
rect 204536 4004 204588 4010
rect 204536 3946 204588 3952
rect 204352 3936 204404 3942
rect 204352 3878 204404 3884
rect 205100 480 205128 6190
rect 205652 4078 205680 104042
rect 205744 9042 205772 110078
rect 206020 99374 206048 110078
rect 206480 104106 206508 110078
rect 207020 104168 207072 104174
rect 207020 104110 207072 104116
rect 206468 104100 206520 104106
rect 206468 104042 206520 104048
rect 205836 99346 206048 99374
rect 205836 69698 205864 99346
rect 205824 69692 205876 69698
rect 205824 69634 205876 69640
rect 205824 44872 205876 44878
rect 205824 44814 205876 44820
rect 205836 16574 205864 44814
rect 205836 16546 206232 16574
rect 205732 9036 205784 9042
rect 205732 8978 205784 8984
rect 205640 4072 205692 4078
rect 205640 4014 205692 4020
rect 206204 480 206232 16546
rect 207032 4146 207060 104110
rect 207124 10334 207152 110078
rect 207308 99374 207336 110078
rect 207676 104174 207704 110078
rect 208412 109034 208440 110092
rect 208320 109006 208440 109034
rect 208504 110078 208794 110106
rect 208872 110078 209254 110106
rect 207664 104168 207716 104174
rect 207664 104110 207716 104116
rect 208320 102814 208348 109006
rect 208308 102808 208360 102814
rect 208308 102750 208360 102756
rect 207216 99346 207336 99374
rect 207216 72486 207244 99346
rect 208504 90370 208532 110078
rect 208872 99374 208900 110078
rect 209608 108662 209636 110092
rect 209884 110078 210082 110106
rect 210160 110078 210450 110106
rect 210528 110078 210818 110106
rect 211278 110078 211476 110106
rect 209596 108656 209648 108662
rect 209596 108598 209648 108604
rect 209780 104168 209832 104174
rect 209780 104110 209832 104116
rect 208596 99346 208900 99374
rect 208492 90364 208544 90370
rect 208492 90306 208544 90312
rect 208596 73846 208624 99346
rect 208584 73840 208636 73846
rect 208584 73782 208636 73788
rect 207204 72480 207256 72486
rect 207204 72422 207256 72428
rect 207112 10328 207164 10334
rect 207112 10270 207164 10276
rect 208584 9036 208636 9042
rect 208584 8978 208636 8984
rect 207388 6316 207440 6322
rect 207388 6258 207440 6264
rect 207020 4140 207072 4146
rect 207020 4082 207072 4088
rect 207400 480 207428 6258
rect 208596 480 208624 8978
rect 209792 6914 209820 104110
rect 209884 10402 209912 110078
rect 210160 99374 210188 110078
rect 210528 104174 210556 110078
rect 211448 104378 211476 110078
rect 211540 110078 211646 110106
rect 211436 104372 211488 104378
rect 211436 104314 211488 104320
rect 210516 104168 210568 104174
rect 210516 104110 210568 104116
rect 211252 104168 211304 104174
rect 211252 104110 211304 104116
rect 209976 99346 210188 99374
rect 209976 75206 210004 99346
rect 209964 75200 210016 75206
rect 209964 75142 210016 75148
rect 211264 49026 211292 104110
rect 211540 101402 211568 110078
rect 211804 107704 211856 107710
rect 211804 107646 211856 107652
rect 211620 104372 211672 104378
rect 211620 104314 211672 104320
rect 211356 101374 211568 101402
rect 211356 82142 211384 101374
rect 211632 96614 211660 104314
rect 211448 96586 211660 96614
rect 211344 82136 211396 82142
rect 211344 82078 211396 82084
rect 211252 49020 211304 49026
rect 211252 48962 211304 48968
rect 209964 47660 210016 47666
rect 209964 47602 210016 47608
rect 209872 10396 209924 10402
rect 209872 10338 209924 10344
rect 209792 6886 209912 6914
rect 209884 5098 209912 6886
rect 209872 5092 209924 5098
rect 209872 5034 209924 5040
rect 209976 3482 210004 47602
rect 211448 21418 211476 96586
rect 211816 29646 211844 107646
rect 212092 104106 212120 110092
rect 212184 110078 212474 110106
rect 212184 104174 212212 110078
rect 212828 107710 212856 110092
rect 212920 110078 213302 110106
rect 213380 110078 213670 110106
rect 212816 107704 212868 107710
rect 212816 107646 212868 107652
rect 212920 105602 212948 110078
rect 213380 109034 213408 110078
rect 213104 109006 213408 109034
rect 212908 105596 212960 105602
rect 212908 105538 212960 105544
rect 212172 104168 212224 104174
rect 212172 104110 212224 104116
rect 212080 104100 212132 104106
rect 212080 104042 212132 104048
rect 213104 99374 213132 109006
rect 214116 107710 214144 110092
rect 214208 110078 214498 110106
rect 214576 110078 214866 110106
rect 215326 110078 215432 110106
rect 213184 107704 213236 107710
rect 213184 107646 213236 107652
rect 214104 107704 214156 107710
rect 214104 107646 214156 107652
rect 212736 99346 213132 99374
rect 212736 89010 212764 99346
rect 212724 89004 212776 89010
rect 212724 88946 212776 88952
rect 213196 76566 213224 107646
rect 214012 104168 214064 104174
rect 214012 104110 214064 104116
rect 214024 80714 214052 104110
rect 214208 99374 214236 110078
rect 214576 104174 214604 110078
rect 214656 107704 214708 107710
rect 214656 107646 214708 107652
rect 214564 104168 214616 104174
rect 214564 104110 214616 104116
rect 214668 99374 214696 107646
rect 215404 107166 215432 110078
rect 215392 107160 215444 107166
rect 215392 107102 215444 107108
rect 215392 106820 215444 106826
rect 215392 106762 215444 106768
rect 214116 99346 214236 99374
rect 214576 99346 214696 99374
rect 214012 80708 214064 80714
rect 214012 80650 214064 80656
rect 213184 76560 213236 76566
rect 213184 76502 213236 76508
rect 211804 29640 211856 29646
rect 211804 29582 211856 29588
rect 211436 21412 211488 21418
rect 211436 21354 211488 21360
rect 214012 21412 214064 21418
rect 214012 21354 214064 21360
rect 210056 20052 210108 20058
rect 210056 19994 210108 20000
rect 210068 16574 210096 19994
rect 210068 16546 211016 16574
rect 209792 3454 210004 3482
rect 209792 480 209820 3454
rect 210988 480 211016 16546
rect 211712 15972 211764 15978
rect 211712 15914 211764 15920
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 15914
rect 213368 7608 213420 7614
rect 213368 7550 213420 7556
rect 213380 480 213408 7550
rect 214024 3482 214052 21354
rect 214116 6186 214144 99346
rect 214576 18630 214604 99346
rect 215404 42090 215432 106762
rect 215496 61402 215524 110214
rect 224960 110162 225012 110168
rect 225144 110220 225446 110226
rect 225196 110214 225446 110220
rect 229126 110214 229416 110242
rect 238956 110226 239246 110242
rect 345216 110226 345506 110242
rect 225144 110162 225196 110168
rect 216140 107710 216168 110092
rect 216232 110078 216522 110106
rect 216784 110078 216890 110106
rect 216968 110078 217350 110106
rect 216128 107704 216180 107710
rect 216128 107646 216180 107652
rect 215576 107160 215628 107166
rect 215576 107102 215628 107108
rect 215484 61396 215536 61402
rect 215484 61338 215536 61344
rect 215392 42084 215444 42090
rect 215392 42026 215444 42032
rect 215392 31136 215444 31142
rect 215392 31078 215444 31084
rect 214564 18624 214616 18630
rect 214564 18566 214616 18572
rect 214104 6180 214156 6186
rect 214104 6122 214156 6128
rect 214024 3454 214512 3482
rect 214484 480 214512 3454
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215404 354 215432 31078
rect 215588 28286 215616 107102
rect 216232 106826 216260 110078
rect 216220 106820 216272 106826
rect 216220 106762 216272 106768
rect 216784 60042 216812 110078
rect 216968 103514 216996 110078
rect 217324 107704 217376 107710
rect 217324 107646 217376 107652
rect 216876 103486 216996 103514
rect 216772 60036 216824 60042
rect 216772 59978 216824 59984
rect 216772 49020 216824 49026
rect 216772 48962 216824 48968
rect 215576 28280 215628 28286
rect 215576 28222 215628 28228
rect 216784 16574 216812 48962
rect 216876 31074 216904 103486
rect 217336 77994 217364 107646
rect 217704 106962 217732 110092
rect 218164 107710 218192 110092
rect 218256 110078 218546 110106
rect 218624 110078 219006 110106
rect 219084 110078 219374 110106
rect 219544 110078 219742 110106
rect 219820 110078 220202 110106
rect 220280 110078 220570 110106
rect 220832 110078 221030 110106
rect 221108 110078 221398 110106
rect 221476 110078 221766 110106
rect 218152 107704 218204 107710
rect 218152 107646 218204 107652
rect 217692 106956 217744 106962
rect 217692 106898 217744 106904
rect 218256 106842 218284 110078
rect 218164 106814 218284 106842
rect 218164 87650 218192 106814
rect 218244 106752 218296 106758
rect 218244 106694 218296 106700
rect 218256 94518 218284 106694
rect 218624 103514 218652 110078
rect 218704 108316 218756 108322
rect 218704 108258 218756 108264
rect 218348 103486 218652 103514
rect 218244 94512 218296 94518
rect 218244 94454 218296 94460
rect 218152 87644 218204 87650
rect 218152 87586 218204 87592
rect 217324 77988 217376 77994
rect 217324 77930 217376 77936
rect 216864 31068 216916 31074
rect 216864 31010 216916 31016
rect 218348 26926 218376 103486
rect 218716 47598 218744 108258
rect 219084 106758 219112 110078
rect 219440 106820 219492 106826
rect 219440 106762 219492 106768
rect 219072 106752 219124 106758
rect 219072 106694 219124 106700
rect 218704 47592 218756 47598
rect 218704 47534 218756 47540
rect 218336 26920 218388 26926
rect 218336 26862 218388 26868
rect 218060 17264 218112 17270
rect 218060 17206 218112 17212
rect 216784 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 3534 218100 17206
rect 219452 7886 219480 106762
rect 219544 11762 219572 110078
rect 219820 103514 219848 110078
rect 220084 107772 220136 107778
rect 220084 107714 220136 107720
rect 219636 103486 219848 103514
rect 219636 98734 219664 103486
rect 219624 98728 219676 98734
rect 219624 98670 219676 98676
rect 220096 57254 220124 107714
rect 220280 106826 220308 110078
rect 220268 106820 220320 106826
rect 220268 106762 220320 106768
rect 220084 57248 220136 57254
rect 220084 57190 220136 57196
rect 219624 51808 219676 51814
rect 219624 51750 219676 51756
rect 219636 16574 219664 51750
rect 219636 16546 220032 16574
rect 219532 11756 219584 11762
rect 219532 11698 219584 11704
rect 219440 7880 219492 7886
rect 219440 7822 219492 7828
rect 218152 5024 218204 5030
rect 218152 4966 218204 4972
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 218164 2530 218192 4966
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 218072 2502 218192 2530
rect 218072 480 218100 2502
rect 219268 480 219296 3470
rect 215638 354 215750 480
rect 215404 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220832 11830 220860 110078
rect 221108 106808 221136 110078
rect 220924 106780 221136 106808
rect 220924 25566 220952 106780
rect 221476 106740 221504 110078
rect 222212 108322 222240 110092
rect 222396 110078 222594 110106
rect 222200 108316 222252 108322
rect 222200 108258 222252 108264
rect 221556 107704 221608 107710
rect 221556 107646 221608 107652
rect 221016 106712 221504 106740
rect 221016 58682 221044 106712
rect 221568 103514 221596 107646
rect 222292 106820 222344 106826
rect 222292 106762 222344 106768
rect 221476 103486 221596 103514
rect 221476 93158 221504 103486
rect 221464 93152 221516 93158
rect 221464 93094 221516 93100
rect 222304 66910 222332 106762
rect 222292 66904 222344 66910
rect 222292 66846 222344 66852
rect 221004 58676 221056 58682
rect 221004 58618 221056 58624
rect 222396 54534 222424 110078
rect 223040 107710 223068 110092
rect 223132 110078 223422 110106
rect 223790 110078 223896 110106
rect 223028 107704 223080 107710
rect 223028 107646 223080 107652
rect 223132 106826 223160 110078
rect 223580 108316 223632 108322
rect 223580 108258 223632 108264
rect 223120 106820 223172 106826
rect 223120 106762 223172 106768
rect 222384 54528 222436 54534
rect 222384 54470 222436 54476
rect 220912 25560 220964 25566
rect 220912 25502 220964 25508
rect 221096 14544 221148 14550
rect 221096 14486 221148 14492
rect 220820 11824 220872 11830
rect 220820 11766 220872 11772
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 14486
rect 222752 7676 222804 7682
rect 222752 7618 222804 7624
rect 222764 480 222792 7618
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 108258
rect 223764 106888 223816 106894
rect 223764 106830 223816 106836
rect 223672 106820 223724 106826
rect 223672 106762 223724 106768
rect 223684 10470 223712 106762
rect 223776 11898 223804 106830
rect 223868 84862 223896 110078
rect 223960 110078 224250 110106
rect 224328 110078 224618 110106
rect 223960 106826 223988 110078
rect 224328 106894 224356 110078
rect 224316 106888 224368 106894
rect 224316 106830 224368 106836
rect 223948 106820 224000 106826
rect 223948 106762 224000 106768
rect 223856 84856 223908 84862
rect 223856 84798 223908 84804
rect 223764 11892 223816 11898
rect 223764 11834 223816 11840
rect 224972 10538 225000 110162
rect 225078 110078 225276 110106
rect 225052 104168 225104 104174
rect 225052 104110 225104 104116
rect 225064 11966 225092 104110
rect 225144 101448 225196 101454
rect 225144 101390 225196 101396
rect 225156 64190 225184 101390
rect 225248 65550 225276 110078
rect 225616 110078 225906 110106
rect 225984 110078 226274 110106
rect 225616 104174 225644 110078
rect 225604 104168 225656 104174
rect 225604 104110 225656 104116
rect 225984 101454 226012 110078
rect 226628 107778 226656 110092
rect 226720 110078 227102 110106
rect 227180 110078 227470 110106
rect 227824 110078 227930 110106
rect 228008 110078 228298 110106
rect 228376 110078 228666 110106
rect 226616 107772 226668 107778
rect 226616 107714 226668 107720
rect 226720 104258 226748 110078
rect 226444 104230 226748 104258
rect 225972 101448 226024 101454
rect 225972 101390 226024 101396
rect 226444 83502 226472 104230
rect 227180 99374 227208 110078
rect 227720 104168 227772 104174
rect 227720 104110 227772 104116
rect 226536 99346 227208 99374
rect 226432 83496 226484 83502
rect 226432 83438 226484 83444
rect 225236 65544 225288 65550
rect 225236 65486 225288 65492
rect 225144 64184 225196 64190
rect 225144 64126 225196 64132
rect 226536 53106 226564 99346
rect 226524 53100 226576 53106
rect 226524 53042 226576 53048
rect 225052 11960 225104 11966
rect 225052 11902 225104 11908
rect 224960 10532 225012 10538
rect 224960 10474 225012 10480
rect 223672 10464 223724 10470
rect 223672 10406 223724 10412
rect 226340 10396 226392 10402
rect 226340 10338 226392 10344
rect 225144 10328 225196 10334
rect 225144 10270 225196 10276
rect 225156 480 225184 10270
rect 226352 480 226380 10338
rect 227536 6180 227588 6186
rect 227536 6122 227588 6128
rect 227548 480 227576 6122
rect 227732 3398 227760 104110
rect 227824 10606 227852 110078
rect 228008 99374 228036 110078
rect 228376 104174 228404 110078
rect 228364 104168 228416 104174
rect 228364 104110 228416 104116
rect 229284 104168 229336 104174
rect 229284 104110 229336 104116
rect 229192 100972 229244 100978
rect 229192 100914 229244 100920
rect 227916 99346 228036 99374
rect 227916 12034 227944 99346
rect 229204 12102 229232 100914
rect 229296 55894 229324 104110
rect 229284 55888 229336 55894
rect 229284 55830 229336 55836
rect 229192 12096 229244 12102
rect 229192 12038 229244 12044
rect 227904 12028 227956 12034
rect 227904 11970 227956 11976
rect 228272 11756 228324 11762
rect 228272 11698 228324 11704
rect 227812 10600 227864 10606
rect 227812 10542 227864 10548
rect 227720 3392 227772 3398
rect 227720 3334 227772 3340
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 11698
rect 229388 10674 229416 110214
rect 238760 110220 238812 110226
rect 238760 110162 238812 110168
rect 238944 110220 239246 110226
rect 238996 110214 239246 110220
rect 345020 110220 345072 110226
rect 238944 110162 238996 110168
rect 345020 110162 345072 110168
rect 345204 110220 345506 110226
rect 345256 110214 345506 110220
rect 345204 110162 345256 110168
rect 229480 100978 229508 110092
rect 229940 108458 229968 110092
rect 230032 110078 230322 110106
rect 229928 108452 229980 108458
rect 229928 108394 229980 108400
rect 230032 104174 230060 110078
rect 230676 109034 230704 110092
rect 230584 109006 230704 109034
rect 230768 110078 231150 110106
rect 231228 110078 231518 110106
rect 231978 110078 232176 110106
rect 230584 106274 230612 109006
rect 230768 106274 230796 110078
rect 230400 106246 230612 106274
rect 230676 106246 230796 106274
rect 230020 104168 230072 104174
rect 230020 104110 230072 104116
rect 230400 101454 230428 106246
rect 230676 101538 230704 106246
rect 230492 101510 230704 101538
rect 230388 101448 230440 101454
rect 230388 101390 230440 101396
rect 229468 100972 229520 100978
rect 229468 100914 229520 100920
rect 229376 10668 229428 10674
rect 229376 10610 229428 10616
rect 229836 7744 229888 7750
rect 229836 7686 229888 7692
rect 229848 480 229876 7686
rect 230492 3330 230520 101510
rect 230572 101448 230624 101454
rect 230572 101390 230624 101396
rect 230584 13190 230612 101390
rect 231228 99374 231256 110078
rect 232044 104168 232096 104174
rect 232044 104110 232096 104116
rect 231952 104100 232004 104106
rect 231952 104042 232004 104048
rect 230676 99346 231256 99374
rect 230676 86290 230704 99346
rect 230664 86284 230716 86290
rect 230664 86226 230716 86232
rect 231964 13326 231992 104042
rect 232056 35222 232084 104110
rect 232044 35216 232096 35222
rect 232044 35158 232096 35164
rect 231952 13320 232004 13326
rect 231952 13262 232004 13268
rect 232148 13258 232176 110078
rect 232332 108526 232360 110092
rect 232424 110078 232714 110106
rect 232792 110078 233174 110106
rect 233252 110078 233542 110106
rect 233620 110078 234002 110106
rect 234080 110078 234370 110106
rect 232320 108520 232372 108526
rect 232320 108462 232372 108468
rect 232424 104174 232452 110078
rect 232412 104168 232464 104174
rect 232412 104110 232464 104116
rect 232792 104106 232820 110078
rect 232780 104100 232832 104106
rect 232780 104042 232832 104048
rect 232136 13252 232188 13258
rect 232136 13194 232188 13200
rect 230572 13184 230624 13190
rect 230572 13126 230624 13132
rect 232044 13116 232096 13122
rect 232044 13058 232096 13064
rect 231032 3460 231084 3466
rect 231032 3402 231084 3408
rect 230480 3324 230532 3330
rect 230480 3266 230532 3272
rect 231044 480 231072 3402
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232056 354 232084 13058
rect 233252 3262 233280 110078
rect 233332 104168 233384 104174
rect 233332 104110 233384 104116
rect 233344 13394 233372 104110
rect 233620 99374 233648 110078
rect 234080 104174 234108 110078
rect 234816 108594 234844 110092
rect 234908 110078 235198 110106
rect 235276 110078 235566 110106
rect 234804 108588 234856 108594
rect 234804 108530 234856 108536
rect 234908 107030 234936 110078
rect 235276 109034 235304 110078
rect 235184 109006 235304 109034
rect 234896 107024 234948 107030
rect 234896 106966 234948 106972
rect 234068 104168 234120 104174
rect 234068 104110 234120 104116
rect 235184 99374 235212 109006
rect 235356 108520 235408 108526
rect 235356 108462 235408 108468
rect 235264 108384 235316 108390
rect 235264 108326 235316 108332
rect 233436 99346 233648 99374
rect 234724 99346 235212 99374
rect 233436 51746 233464 99346
rect 234724 82210 234752 99346
rect 234712 82204 234764 82210
rect 234712 82146 234764 82152
rect 233424 51740 233476 51746
rect 233424 51682 233476 51688
rect 233424 35216 233476 35222
rect 233424 35158 233476 35164
rect 233332 13388 233384 13394
rect 233332 13330 233384 13336
rect 233240 3256 233292 3262
rect 233240 3198 233292 3204
rect 233436 480 233464 35158
rect 235276 5030 235304 108326
rect 235368 14482 235396 108462
rect 235448 107704 235500 107710
rect 235448 107646 235500 107652
rect 235460 94586 235488 107646
rect 236012 106274 236040 110092
rect 236380 107710 236408 110092
rect 236472 110078 236854 110106
rect 236932 110078 237222 110106
rect 237484 110078 237590 110106
rect 237760 110078 238050 110106
rect 236368 107704 236420 107710
rect 236368 107646 236420 107652
rect 236012 106246 236316 106274
rect 236092 99272 236144 99278
rect 236092 99214 236144 99220
rect 236104 96014 236132 99214
rect 236092 96008 236144 96014
rect 236092 95950 236144 95956
rect 235448 94580 235500 94586
rect 235448 94522 235500 94528
rect 236288 39370 236316 106246
rect 236472 99278 236500 110078
rect 236644 107704 236696 107710
rect 236644 107646 236696 107652
rect 236460 99272 236512 99278
rect 236460 99214 236512 99220
rect 236656 65618 236684 107646
rect 236932 101522 236960 110078
rect 236920 101516 236972 101522
rect 236920 101458 236972 101464
rect 237484 93226 237512 110078
rect 237760 99374 237788 110078
rect 238116 107840 238168 107846
rect 238116 107782 238168 107788
rect 238024 107772 238076 107778
rect 238024 107714 238076 107720
rect 237576 99346 237788 99374
rect 237472 93220 237524 93226
rect 237472 93162 237524 93168
rect 237576 76634 237604 99346
rect 237564 76628 237616 76634
rect 237564 76570 237616 76576
rect 236644 65612 236696 65618
rect 236644 65554 236696 65560
rect 236276 39364 236328 39370
rect 236276 39306 236328 39312
rect 236000 36644 236052 36650
rect 236000 36586 236052 36592
rect 236012 16574 236040 36586
rect 238036 36582 238064 107714
rect 238128 89078 238156 107782
rect 238404 107710 238432 110092
rect 238392 107704 238444 107710
rect 238392 107646 238444 107652
rect 238116 89072 238168 89078
rect 238116 89014 238168 89020
rect 238772 37942 238800 110162
rect 238878 110078 239076 110106
rect 238852 104168 238904 104174
rect 238852 104110 238904 104116
rect 238864 64258 238892 104110
rect 238944 100768 238996 100774
rect 238944 100710 238996 100716
rect 238956 90438 238984 100710
rect 239048 91866 239076 110078
rect 239324 110078 239614 110106
rect 239784 110078 240074 110106
rect 239324 104174 239352 110078
rect 239312 104168 239364 104174
rect 239312 104110 239364 104116
rect 239784 100774 239812 110078
rect 240428 107778 240456 110092
rect 240520 110078 240902 110106
rect 240416 107772 240468 107778
rect 240416 107714 240468 107720
rect 239772 100768 239824 100774
rect 239772 100710 239824 100716
rect 240520 99374 240548 110078
rect 241256 107846 241284 110092
rect 241532 110078 241638 110106
rect 241716 110078 242098 110106
rect 242176 110078 242466 110106
rect 242926 110078 243124 110106
rect 241244 107840 241296 107846
rect 241244 107782 241296 107788
rect 240244 99346 240548 99374
rect 240244 97374 240272 99346
rect 240232 97368 240284 97374
rect 240232 97310 240284 97316
rect 239036 91860 239088 91866
rect 239036 91802 239088 91808
rect 238944 90432 238996 90438
rect 238944 90374 238996 90380
rect 238852 64252 238904 64258
rect 238852 64194 238904 64200
rect 241532 46238 241560 110078
rect 241716 109034 241744 110078
rect 242176 109034 242204 110078
rect 241624 109006 241744 109034
rect 241992 109006 242204 109034
rect 241624 50386 241652 109006
rect 241992 99374 242020 109006
rect 242164 107704 242216 107710
rect 242164 107646 242216 107652
rect 241716 99346 242020 99374
rect 241716 87718 241744 99346
rect 241704 87712 241756 87718
rect 241704 87654 241756 87660
rect 242176 83570 242204 107646
rect 243096 104650 243124 110078
rect 243188 110078 243294 110106
rect 243464 110078 243754 110106
rect 243832 110078 244122 110106
rect 244384 110078 244490 110106
rect 243084 104644 243136 104650
rect 243084 104586 243136 104592
rect 243084 104440 243136 104446
rect 243084 104382 243136 104388
rect 242992 104168 243044 104174
rect 242992 104110 243044 104116
rect 242900 101448 242952 101454
rect 242900 101390 242952 101396
rect 242164 83564 242216 83570
rect 242164 83506 242216 83512
rect 242912 53174 242940 101390
rect 243004 73914 243032 104110
rect 243096 75274 243124 104382
rect 243188 101454 243216 110078
rect 243176 101448 243228 101454
rect 243176 101390 243228 101396
rect 243464 99374 243492 110078
rect 243832 104174 243860 110078
rect 243820 104168 243872 104174
rect 243820 104110 243872 104116
rect 244384 100094 244412 110078
rect 244936 107710 244964 110092
rect 245028 110078 245318 110106
rect 245778 110078 245884 110106
rect 244924 107704 244976 107710
rect 244924 107646 244976 107652
rect 245028 103514 245056 110078
rect 245752 106820 245804 106826
rect 245752 106762 245804 106768
rect 244476 103486 245056 103514
rect 244372 100088 244424 100094
rect 244372 100030 244424 100036
rect 243188 99346 243492 99374
rect 243188 86358 243216 99346
rect 243176 86352 243228 86358
rect 243176 86294 243228 86300
rect 243084 75268 243136 75274
rect 243084 75210 243136 75216
rect 242992 73908 243044 73914
rect 242992 73850 243044 73856
rect 244476 72554 244504 103486
rect 244464 72548 244516 72554
rect 244464 72490 244516 72496
rect 245764 54602 245792 106762
rect 245856 62898 245884 110078
rect 246132 107098 246160 110092
rect 246224 110078 246514 110106
rect 246592 110078 246974 110106
rect 246120 107092 246172 107098
rect 246120 107034 246172 107040
rect 246224 103514 246252 110078
rect 246592 106826 246620 110078
rect 247224 108180 247276 108186
rect 247224 108122 247276 108128
rect 246580 106820 246632 106826
rect 246580 106762 246632 106768
rect 247132 106820 247184 106826
rect 247132 106762 247184 106768
rect 247040 104168 247092 104174
rect 247040 104110 247092 104116
rect 245948 103486 246252 103514
rect 245844 62892 245896 62898
rect 245844 62834 245896 62840
rect 245752 54596 245804 54602
rect 245752 54538 245804 54544
rect 242900 53168 242952 53174
rect 242900 53110 242952 53116
rect 241612 50380 241664 50386
rect 241612 50322 241664 50328
rect 241520 46232 241572 46238
rect 241520 46174 241572 46180
rect 245948 40730 245976 103486
rect 245936 40724 245988 40730
rect 245936 40666 245988 40672
rect 242900 39364 242952 39370
rect 242900 39306 242952 39312
rect 238760 37936 238812 37942
rect 238760 37878 238812 37884
rect 238024 36576 238076 36582
rect 238024 36518 238076 36524
rect 236012 16546 236592 16574
rect 235356 14476 235408 14482
rect 235356 14418 235408 14424
rect 235264 5024 235316 5030
rect 235264 4966 235316 4972
rect 235816 4956 235868 4962
rect 235816 4898 235868 4904
rect 234620 3188 234672 3194
rect 234620 3130 234672 3136
rect 234632 480 234660 3130
rect 235828 480 235856 4898
rect 232198 354 232310 480
rect 232056 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 240140 11824 240192 11830
rect 240140 11766 240192 11772
rect 239312 9104 239364 9110
rect 239312 9046 239364 9052
rect 238116 3596 238168 3602
rect 238116 3538 238168 3544
rect 238128 480 238156 3538
rect 239324 480 239352 9046
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 11766
rect 241704 3664 241756 3670
rect 241704 3606 241756 3612
rect 241716 480 241744 3606
rect 242912 3534 242940 39306
rect 247052 16574 247080 104110
rect 247144 69766 247172 106762
rect 247236 104242 247264 108122
rect 247328 105670 247356 110092
rect 247512 110078 247802 110106
rect 247880 110078 248170 110106
rect 247316 105664 247368 105670
rect 247316 105606 247368 105612
rect 247224 104236 247276 104242
rect 247224 104178 247276 104184
rect 247512 103514 247540 110078
rect 247684 108452 247736 108458
rect 247684 108394 247736 108400
rect 247236 103486 247540 103514
rect 247236 80782 247264 103486
rect 247224 80776 247276 80782
rect 247224 80718 247276 80724
rect 247132 69760 247184 69766
rect 247132 69702 247184 69708
rect 247052 16546 247632 16574
rect 246396 6452 246448 6458
rect 246396 6394 246448 6400
rect 242992 6384 243044 6390
rect 242992 6326 243044 6332
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 243004 3210 243032 6326
rect 245200 3732 245252 3738
rect 245200 3674 245252 3680
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242912 3182 243032 3210
rect 242912 480 242940 3182
rect 244108 480 244136 3470
rect 245212 480 245240 3674
rect 246408 480 246436 6394
rect 247604 480 247632 16546
rect 247696 6322 247724 108394
rect 247880 106826 247908 110078
rect 248524 108186 248552 110092
rect 248616 110078 248998 110106
rect 249076 110078 249366 110106
rect 248512 108180 248564 108186
rect 248512 108122 248564 108128
rect 248616 106842 248644 110078
rect 247868 106820 247920 106826
rect 247868 106762 247920 106768
rect 248524 106814 248644 106842
rect 248524 79422 248552 106814
rect 249076 103514 249104 110078
rect 249812 108526 249840 110092
rect 249996 110078 250194 110106
rect 249800 108520 249852 108526
rect 249800 108462 249852 108468
rect 249892 106820 249944 106826
rect 249892 106762 249944 106768
rect 248616 103486 249104 103514
rect 248512 79416 248564 79422
rect 248512 79358 248564 79364
rect 248616 68406 248644 103486
rect 249904 102882 249932 106762
rect 249892 102876 249944 102882
rect 249892 102818 249944 102824
rect 248604 68400 248656 68406
rect 248604 68342 248656 68348
rect 249996 22778 250024 110078
rect 250444 108520 250496 108526
rect 250444 108462 250496 108468
rect 249984 22772 250036 22778
rect 249984 22714 250036 22720
rect 250456 20058 250484 108462
rect 250536 107704 250588 107710
rect 250536 107646 250588 107652
rect 250548 100162 250576 107646
rect 250640 105738 250668 110092
rect 250732 110078 251022 110106
rect 251284 110078 251390 110106
rect 250732 106826 250760 110078
rect 250720 106820 250772 106826
rect 250720 106762 250772 106768
rect 250628 105732 250680 105738
rect 250628 105674 250680 105680
rect 251180 101448 251232 101454
rect 251180 101390 251232 101396
rect 250536 100156 250588 100162
rect 250536 100098 250588 100104
rect 250444 20052 250496 20058
rect 250444 19994 250496 20000
rect 247684 6316 247736 6322
rect 247684 6258 247736 6264
rect 249984 5024 250036 5030
rect 249984 4966 250036 4972
rect 248788 3800 248840 3806
rect 248788 3742 248840 3748
rect 248800 480 248828 3742
rect 249996 480 250024 4966
rect 251192 480 251220 101390
rect 251284 24138 251312 110078
rect 251836 104310 251864 110092
rect 251928 110078 252218 110106
rect 252572 110078 252678 110106
rect 252756 110078 253046 110106
rect 251824 104304 251876 104310
rect 251824 104246 251876 104252
rect 251928 104122 251956 110078
rect 252008 108044 252060 108050
rect 252008 107986 252060 107992
rect 251376 104094 251956 104122
rect 251376 101590 251404 104094
rect 252020 103514 252048 107986
rect 252572 104514 252600 110078
rect 252756 106842 252784 110078
rect 253204 108588 253256 108594
rect 253204 108530 253256 108536
rect 252664 106814 252784 106842
rect 252560 104508 252612 104514
rect 252560 104450 252612 104456
rect 251836 103486 252048 103514
rect 251364 101584 251416 101590
rect 251364 101526 251416 101532
rect 251272 24132 251324 24138
rect 251272 24074 251324 24080
rect 251836 15910 251864 103486
rect 252664 42158 252692 106814
rect 252744 106752 252796 106758
rect 252744 106694 252796 106700
rect 252756 84930 252784 106694
rect 252836 104508 252888 104514
rect 252836 104450 252888 104456
rect 252744 84924 252796 84930
rect 252744 84866 252796 84872
rect 252652 42152 252704 42158
rect 252652 42094 252704 42100
rect 252848 25634 252876 104450
rect 252836 25628 252888 25634
rect 252836 25570 252888 25576
rect 252560 22772 252612 22778
rect 252560 22714 252612 22720
rect 252572 16574 252600 22714
rect 252572 16546 253152 16574
rect 251824 15904 251876 15910
rect 251824 15846 251876 15852
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 252388 480 252416 3810
rect 253124 3482 253152 16546
rect 253216 6254 253244 108530
rect 253400 107710 253428 110092
rect 253584 110078 253874 110106
rect 254044 110078 254242 110106
rect 254320 110078 254702 110106
rect 254780 110078 255070 110106
rect 253388 107704 253440 107710
rect 253388 107646 253440 107652
rect 253584 106758 253612 110078
rect 253940 106820 253992 106826
rect 253940 106762 253992 106768
rect 253572 106752 253624 106758
rect 253572 106694 253624 106700
rect 253952 78062 253980 106762
rect 253940 78056 253992 78062
rect 253940 77998 253992 78004
rect 254044 66978 254072 110078
rect 254320 103514 254348 110078
rect 254780 106826 254808 110078
rect 254768 106820 254820 106826
rect 254768 106762 254820 106768
rect 255320 106820 255372 106826
rect 255320 106762 255372 106768
rect 254136 103486 254348 103514
rect 254136 98802 254164 103486
rect 254124 98796 254176 98802
rect 254124 98738 254176 98744
rect 254124 78192 254176 78198
rect 254124 78134 254176 78140
rect 254032 66972 254084 66978
rect 254032 66914 254084 66920
rect 254136 16574 254164 78134
rect 255332 26994 255360 106762
rect 255424 71058 255452 110092
rect 255516 110078 255898 110106
rect 255976 110078 256266 110106
rect 256726 110078 257016 110106
rect 255516 97442 255544 110078
rect 255976 106826 256004 110078
rect 256056 107704 256108 107710
rect 256056 107646 256108 107652
rect 255964 106820 256016 106826
rect 255964 106762 256016 106768
rect 256068 103514 256096 107646
rect 256884 106888 256936 106894
rect 256884 106830 256936 106836
rect 256792 106820 256844 106826
rect 256792 106762 256844 106768
rect 255976 103486 256096 103514
rect 255504 97436 255556 97442
rect 255504 97378 255556 97384
rect 255412 71052 255464 71058
rect 255412 70994 255464 71000
rect 255976 32434 256004 103486
rect 255964 32428 256016 32434
rect 255964 32370 256016 32376
rect 256804 28354 256832 106762
rect 256792 28348 256844 28354
rect 256792 28290 256844 28296
rect 255320 26988 255372 26994
rect 255320 26930 255372 26936
rect 256896 19990 256924 106830
rect 256988 102950 257016 110078
rect 257080 107710 257108 110092
rect 257172 110078 257462 110106
rect 257632 110078 257922 110106
rect 257068 107704 257120 107710
rect 257068 107646 257120 107652
rect 257172 106826 257200 110078
rect 257436 108180 257488 108186
rect 257436 108122 257488 108128
rect 257344 108112 257396 108118
rect 257344 108054 257396 108060
rect 257160 106820 257212 106826
rect 257160 106762 257212 106768
rect 256976 102944 257028 102950
rect 256976 102886 257028 102892
rect 256884 19984 256936 19990
rect 256884 19926 256936 19932
rect 254136 16546 254256 16574
rect 253204 6248 253256 6254
rect 253204 6190 253256 6196
rect 253124 3454 253520 3482
rect 253492 480 253520 3454
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 256700 15904 256752 15910
rect 256700 15846 256752 15852
rect 255872 3936 255924 3942
rect 255872 3878 255924 3884
rect 255884 480 255912 3878
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 15846
rect 257356 4826 257384 108054
rect 257448 96082 257476 108122
rect 257632 106894 257660 110078
rect 258276 108186 258304 110092
rect 258368 110078 258750 110106
rect 258264 108180 258316 108186
rect 258264 108122 258316 108128
rect 257620 106888 257672 106894
rect 257620 106830 257672 106836
rect 258368 103514 258396 110078
rect 259104 108118 259132 110092
rect 259092 108112 259144 108118
rect 259092 108054 259144 108060
rect 259564 108050 259592 110092
rect 259656 110078 259946 110106
rect 260024 110078 260314 110106
rect 260392 110078 260774 110106
rect 260852 110078 261142 110106
rect 261220 110078 261602 110106
rect 261680 110078 261970 110106
rect 259552 108044 259604 108050
rect 259552 107986 259604 107992
rect 259460 106956 259512 106962
rect 259460 106898 259512 106904
rect 258184 103486 258396 103514
rect 257436 96076 257488 96082
rect 257436 96018 257488 96024
rect 258184 29714 258212 103486
rect 258172 29708 258224 29714
rect 258172 29650 258224 29656
rect 258080 25560 258132 25566
rect 258080 25502 258132 25508
rect 258092 16574 258120 25502
rect 258092 16546 258304 16574
rect 257344 4820 257396 4826
rect 257344 4762 257396 4768
rect 258276 480 258304 16546
rect 259472 3534 259500 106898
rect 259552 106820 259604 106826
rect 259552 106762 259604 106768
rect 259564 17338 259592 106762
rect 259656 33794 259684 110078
rect 260024 103514 260052 110078
rect 260392 106826 260420 110078
rect 260380 106820 260432 106826
rect 260380 106762 260432 106768
rect 259748 103486 260052 103514
rect 259748 43518 259776 103486
rect 259736 43512 259788 43518
rect 259736 43454 259788 43460
rect 259644 33788 259696 33794
rect 259644 33730 259696 33736
rect 259552 17332 259604 17338
rect 259552 17274 259604 17280
rect 260852 4894 260880 110078
rect 261220 106842 261248 110078
rect 260944 106814 261248 106842
rect 260944 8974 260972 106814
rect 261680 103514 261708 110078
rect 262324 108594 262352 110092
rect 262416 110078 262798 110106
rect 262312 108588 262364 108594
rect 262312 108530 262364 108536
rect 262416 103514 262444 110078
rect 263152 108458 263180 110092
rect 263626 110078 263916 110106
rect 263140 108452 263192 108458
rect 263140 108394 263192 108400
rect 263888 104378 263916 110078
rect 263876 104372 263928 104378
rect 263876 104314 263928 104320
rect 263692 104236 263744 104242
rect 263692 104178 263744 104184
rect 261036 103486 261708 103514
rect 262324 103486 262444 103514
rect 261036 18698 261064 103486
rect 262324 44878 262352 103486
rect 262312 44872 262364 44878
rect 262312 44814 262364 44820
rect 261116 24132 261168 24138
rect 261116 24074 261168 24080
rect 261024 18692 261076 18698
rect 261024 18634 261076 18640
rect 261128 16574 261156 24074
rect 261128 16546 261800 16574
rect 260932 8968 260984 8974
rect 260932 8910 260984 8916
rect 260840 4888 260892 4894
rect 260840 4830 260892 4836
rect 259552 4004 259604 4010
rect 259552 3946 259604 3952
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 259564 1986 259592 3946
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 259472 1958 259592 1986
rect 259472 480 259500 1958
rect 260668 480 260696 3470
rect 261772 480 261800 16546
rect 263704 15978 263732 104178
rect 263980 99374 264008 110092
rect 264348 108526 264376 110092
rect 264440 110078 264822 110106
rect 264336 108520 264388 108526
rect 264336 108462 264388 108468
rect 264244 107704 264296 107710
rect 264244 107646 264296 107652
rect 264060 104372 264112 104378
rect 264060 104314 264112 104320
rect 263796 99346 264008 99374
rect 263796 47666 263824 99346
rect 264072 96614 264100 104314
rect 263888 96586 264100 96614
rect 263784 47660 263836 47666
rect 263784 47602 263836 47608
rect 263784 18624 263836 18630
rect 263784 18566 263836 18572
rect 263692 15972 263744 15978
rect 263692 15914 263744 15920
rect 263796 6914 263824 18566
rect 263888 9042 263916 96586
rect 263876 9036 263928 9042
rect 263876 8978 263928 8984
rect 264256 7614 264284 107646
rect 264440 104242 264468 110078
rect 265176 107710 265204 110092
rect 265268 110078 265650 110106
rect 265728 110078 266018 110106
rect 266386 110078 266492 110106
rect 265164 107704 265216 107710
rect 265164 107646 265216 107652
rect 264428 104236 264480 104242
rect 264428 104178 264480 104184
rect 265072 104236 265124 104242
rect 265072 104178 265124 104184
rect 265084 31142 265112 104178
rect 265268 99374 265296 110078
rect 265624 108452 265676 108458
rect 265624 108394 265676 108400
rect 265176 99346 265296 99374
rect 265072 31136 265124 31142
rect 265072 31078 265124 31084
rect 265176 21418 265204 99346
rect 265164 21412 265216 21418
rect 265164 21354 265216 21360
rect 265636 9110 265664 108394
rect 265728 104242 265756 110078
rect 265716 104236 265768 104242
rect 265716 104178 265768 104184
rect 266464 49026 266492 110078
rect 266832 108390 266860 110092
rect 266924 110078 267214 110106
rect 267384 110078 267674 110106
rect 267844 110078 268042 110106
rect 268120 110078 268502 110106
rect 266820 108384 266872 108390
rect 266820 108326 266872 108332
rect 266544 104236 266596 104242
rect 266544 104178 266596 104184
rect 266556 51814 266584 104178
rect 266924 99374 266952 110078
rect 267384 104242 267412 110078
rect 267372 104236 267424 104242
rect 267372 104178 267424 104184
rect 266648 99346 266952 99374
rect 266544 51808 266596 51814
rect 266544 51750 266596 51756
rect 266452 49020 266504 49026
rect 266452 48962 266504 48968
rect 266648 17270 266676 99346
rect 266636 17264 266688 17270
rect 266636 17206 266688 17212
rect 267844 14550 267872 110078
rect 268120 99374 268148 110078
rect 268856 108322 268884 110092
rect 268844 108316 268896 108322
rect 268844 108258 268896 108264
rect 269224 107710 269252 110092
rect 269316 110078 269698 110106
rect 269776 110078 270066 110106
rect 268384 107704 268436 107710
rect 268384 107646 268436 107652
rect 269212 107704 269264 107710
rect 269212 107646 269264 107652
rect 267936 99346 268148 99374
rect 267832 14544 267884 14550
rect 267832 14486 267884 14492
rect 267740 10464 267792 10470
rect 267740 10406 267792 10412
rect 265624 9104 265676 9110
rect 265624 9046 265676 9052
rect 264244 7608 264296 7614
rect 264244 7550 264296 7556
rect 263796 6886 264192 6914
rect 262956 4072 263008 4078
rect 262956 4014 263008 4020
rect 262968 480 262996 4014
rect 264164 480 264192 6886
rect 265348 4140 265400 4146
rect 265348 4082 265400 4088
rect 265360 480 265388 4082
rect 266544 3392 266596 3398
rect 266544 3334 266596 3340
rect 266556 480 266584 3334
rect 267752 480 267780 10406
rect 267936 7682 267964 99346
rect 268396 10334 268424 107646
rect 269316 104258 269344 110078
rect 269776 109034 269804 110078
rect 269224 104230 269344 104258
rect 269684 109006 269804 109034
rect 269224 10402 269252 104230
rect 269684 99374 269712 109006
rect 270512 107710 270540 110092
rect 270604 110078 270894 110106
rect 270972 110078 271262 110106
rect 271432 110078 271722 110106
rect 269764 107704 269816 107710
rect 269764 107646 269816 107652
rect 270500 107704 270552 107710
rect 270500 107646 270552 107652
rect 269316 99346 269712 99374
rect 269212 10396 269264 10402
rect 269212 10338 269264 10344
rect 268384 10328 268436 10334
rect 268384 10270 268436 10276
rect 267924 7676 267976 7682
rect 267924 7618 267976 7624
rect 269316 6186 269344 99346
rect 269776 11762 269804 107646
rect 269764 11756 269816 11762
rect 269764 11698 269816 11704
rect 270604 7750 270632 110078
rect 270684 104236 270736 104242
rect 270684 104178 270736 104184
rect 270696 13122 270724 104178
rect 270972 99374 271000 110078
rect 271144 107704 271196 107710
rect 271144 107646 271196 107652
rect 270880 99346 271000 99374
rect 270684 13116 270736 13122
rect 270684 13058 270736 13064
rect 270776 13116 270828 13122
rect 270776 13058 270828 13064
rect 270592 7744 270644 7750
rect 270592 7686 270644 7692
rect 269304 6180 269356 6186
rect 269304 6122 269356 6128
rect 268844 3324 268896 3330
rect 268844 3266 268896 3272
rect 268856 480 268884 3266
rect 270040 3256 270092 3262
rect 270040 3198 270092 3204
rect 270052 480 270080 3198
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 13058
rect 270880 3466 270908 99346
rect 271156 35222 271184 107646
rect 271432 104242 271460 110078
rect 272076 107710 272104 110092
rect 272168 110078 272550 110106
rect 272628 110078 272918 110106
rect 273286 110078 273484 110106
rect 272064 107704 272116 107710
rect 272064 107646 272116 107652
rect 271420 104236 271472 104242
rect 271420 104178 271472 104184
rect 271972 104236 272024 104242
rect 271972 104178 272024 104184
rect 271144 35216 271196 35222
rect 271144 35158 271196 35164
rect 271984 4962 272012 104178
rect 272168 99374 272196 110078
rect 272628 104242 272656 110078
rect 273352 106820 273404 106826
rect 273352 106762 273404 106768
rect 272616 104236 272668 104242
rect 272616 104178 272668 104184
rect 272076 99346 272196 99374
rect 271972 4956 272024 4962
rect 271972 4898 272024 4904
rect 270868 3460 270920 3466
rect 270868 3402 270920 3408
rect 272076 3194 272104 99346
rect 273364 11830 273392 106762
rect 273456 36650 273484 110078
rect 273548 110078 273746 110106
rect 273824 110078 274114 110106
rect 274192 110078 274574 110106
rect 274744 110078 274942 110106
rect 275020 110078 275310 110106
rect 275388 110078 275770 110106
rect 276032 110078 276138 110106
rect 276216 110078 276598 110106
rect 273444 36644 273496 36650
rect 273444 36586 273496 36592
rect 273352 11824 273404 11830
rect 273352 11766 273404 11772
rect 273548 3602 273576 110078
rect 273824 108458 273852 110078
rect 273812 108452 273864 108458
rect 273812 108394 273864 108400
rect 273904 108452 273956 108458
rect 273904 108394 273956 108400
rect 273916 15910 273944 108394
rect 274192 106826 274220 110078
rect 274640 108316 274692 108322
rect 274640 108258 274692 108264
rect 274180 106820 274232 106826
rect 274180 106762 274232 106768
rect 273904 15904 273956 15910
rect 273904 15846 273956 15852
rect 273536 3596 273588 3602
rect 273536 3538 273588 3544
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 274652 3482 274680 108258
rect 274744 3670 274772 110078
rect 275020 106842 275048 110078
rect 274836 106814 275048 106842
rect 274836 16574 274864 106814
rect 275388 103514 275416 110078
rect 276032 103562 276060 110078
rect 276216 106978 276244 110078
rect 276124 106950 276244 106978
rect 274928 103486 275416 103514
rect 276020 103556 276072 103562
rect 276020 103498 276072 103504
rect 274928 39370 274956 103486
rect 274916 39364 274968 39370
rect 274916 39306 274968 39312
rect 274836 16546 274956 16574
rect 274928 6390 274956 16546
rect 276124 6458 276152 106950
rect 276952 104174 276980 110092
rect 277426 110078 277532 110106
rect 277400 104236 277452 104242
rect 277400 104178 277452 104184
rect 276940 104168 276992 104174
rect 276940 104110 276992 104116
rect 276204 103556 276256 103562
rect 276204 103498 276256 103504
rect 276112 6452 276164 6458
rect 276112 6394 276164 6400
rect 274916 6384 274968 6390
rect 274916 6326 274968 6332
rect 276216 3738 276244 103498
rect 277412 101454 277440 104178
rect 277400 101448 277452 101454
rect 277400 101390 277452 101396
rect 277504 3806 277532 110078
rect 277688 110078 277794 110106
rect 277872 110078 278162 110106
rect 278240 110078 278622 110106
rect 277584 106820 277636 106826
rect 277584 106762 277636 106768
rect 277596 3874 277624 106762
rect 277688 5030 277716 110078
rect 277768 108384 277820 108390
rect 277768 108326 277820 108332
rect 277780 16574 277808 108326
rect 277872 104242 277900 110078
rect 278240 106826 278268 110078
rect 278780 108520 278832 108526
rect 278780 108462 278832 108468
rect 278228 106820 278280 106826
rect 278228 106762 278280 106768
rect 277860 104236 277912 104242
rect 277860 104178 277912 104184
rect 277780 16546 278360 16574
rect 277676 5024 277728 5030
rect 277676 4966 277728 4972
rect 277584 3868 277636 3874
rect 277584 3810 277636 3816
rect 277492 3800 277544 3806
rect 277492 3742 277544 3748
rect 276204 3732 276256 3738
rect 276204 3674 276256 3680
rect 274732 3664 274784 3670
rect 274732 3606 274784 3612
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 272064 3188 272116 3194
rect 272064 3130 272116 3136
rect 272444 480 272472 3470
rect 273628 3460 273680 3466
rect 274652 3454 274864 3482
rect 273628 3402 273680 3408
rect 273640 480 273668 3402
rect 274836 480 274864 3454
rect 276032 480 276060 3606
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 277136 480 277164 3538
rect 278332 480 278360 16546
rect 278792 490 278820 108462
rect 278872 106820 278924 106826
rect 278872 106762 278924 106768
rect 278884 3942 278912 106762
rect 278976 22778 279004 110092
rect 279068 110078 279450 110106
rect 279528 110078 279818 110106
rect 279068 78198 279096 110078
rect 279528 106826 279556 110078
rect 280172 108458 280200 110092
rect 280264 110078 280646 110106
rect 280724 110078 281014 110106
rect 280160 108452 280212 108458
rect 280160 108394 280212 108400
rect 279516 106820 279568 106826
rect 279516 106762 279568 106768
rect 279056 78192 279108 78198
rect 279056 78134 279108 78140
rect 280264 25566 280292 110078
rect 280724 103514 280752 110078
rect 281460 106962 281488 110092
rect 281540 108452 281592 108458
rect 281540 108394 281592 108400
rect 281448 106956 281500 106962
rect 281448 106898 281500 106904
rect 280356 103486 280752 103514
rect 280252 25560 280304 25566
rect 280252 25502 280304 25508
rect 278964 22772 279016 22778
rect 278964 22714 279016 22720
rect 280356 4010 280384 103486
rect 280344 4004 280396 4010
rect 280344 3946 280396 3952
rect 280712 4004 280764 4010
rect 280712 3946 280764 3952
rect 278872 3936 278924 3942
rect 278872 3878 278924 3884
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278792 462 279096 490
rect 280724 480 280752 3946
rect 279068 354 279096 462
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 108394
rect 281724 106888 281776 106894
rect 281724 106830 281776 106836
rect 281632 106820 281684 106826
rect 281632 106762 281684 106768
rect 281644 4078 281672 106762
rect 281736 18630 281764 106830
rect 281828 24138 281856 110092
rect 281920 110078 282210 110106
rect 282288 110078 282670 110106
rect 282932 110078 283038 110106
rect 283116 110078 283498 110106
rect 283576 110078 283866 110106
rect 281920 106826 281948 110078
rect 282288 106894 282316 110078
rect 282276 106888 282328 106894
rect 282276 106830 282328 106836
rect 281908 106820 281960 106826
rect 281908 106762 281960 106768
rect 281816 24132 281868 24138
rect 281816 24074 281868 24080
rect 281724 18624 281776 18630
rect 281724 18566 281776 18572
rect 282932 4146 282960 110078
rect 283116 106842 283144 110078
rect 283024 106814 283144 106842
rect 282920 4140 282972 4146
rect 282920 4082 282972 4088
rect 281632 4072 281684 4078
rect 281632 4014 281684 4020
rect 283024 3398 283052 106814
rect 283576 103514 283604 110078
rect 283116 103486 283604 103514
rect 283116 10470 283144 103486
rect 283104 10464 283156 10470
rect 283104 10406 283156 10412
rect 283104 4072 283156 4078
rect 283104 4014 283156 4020
rect 283012 3392 283064 3398
rect 283012 3334 283064 3340
rect 283116 480 283144 4014
rect 284312 3330 284340 110092
rect 284496 110078 284694 110106
rect 284772 110078 285062 110106
rect 285232 110078 285522 110106
rect 285784 110078 285890 110106
rect 284392 106820 284444 106826
rect 284392 106762 284444 106768
rect 284404 3534 284432 106762
rect 284392 3528 284444 3534
rect 284392 3470 284444 3476
rect 284300 3324 284352 3330
rect 284300 3266 284352 3272
rect 284496 3262 284524 110078
rect 284772 103514 284800 110078
rect 285232 106826 285260 110078
rect 285680 108860 285732 108866
rect 285680 108802 285732 108808
rect 285692 108322 285720 108802
rect 285680 108316 285732 108322
rect 285680 108258 285732 108264
rect 285220 106820 285272 106826
rect 285220 106762 285272 106768
rect 284588 103486 284800 103514
rect 284588 13122 284616 103486
rect 284576 13116 284628 13122
rect 284576 13058 284628 13064
rect 285404 4140 285456 4146
rect 285404 4082 285456 4088
rect 284484 3256 284536 3262
rect 284484 3198 284536 3204
rect 284300 3052 284352 3058
rect 284300 2994 284352 3000
rect 284312 480 284340 2994
rect 285416 480 285444 4082
rect 285784 3466 285812 110078
rect 286336 108866 286364 110092
rect 286428 110078 286718 110106
rect 287086 110078 287192 110106
rect 286324 108860 286376 108866
rect 286324 108802 286376 108808
rect 286428 108746 286456 110078
rect 285876 108718 286456 108746
rect 285876 3670 285904 108718
rect 285956 108588 286008 108594
rect 285956 108530 286008 108536
rect 285968 16574 285996 108530
rect 285968 16546 286640 16574
rect 285864 3664 285916 3670
rect 285864 3606 285916 3612
rect 285772 3460 285824 3466
rect 285772 3402 285824 3408
rect 286612 480 286640 16546
rect 287164 3602 287192 110078
rect 287532 108390 287560 110092
rect 287900 108526 287928 110092
rect 287992 110078 288374 110106
rect 287888 108520 287940 108526
rect 287888 108462 287940 108468
rect 287520 108384 287572 108390
rect 287520 108326 287572 108332
rect 287992 107930 288020 110078
rect 288728 108458 288756 110092
rect 288820 110078 289110 110106
rect 289188 110078 289570 110106
rect 288716 108452 288768 108458
rect 288716 108394 288768 108400
rect 287256 107902 288020 107930
rect 287256 4010 287284 107902
rect 287428 107840 287480 107846
rect 287428 107782 287480 107788
rect 287244 4004 287296 4010
rect 287244 3946 287296 3952
rect 287152 3596 287204 3602
rect 287152 3538 287204 3544
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287440 354 287468 107782
rect 288440 107772 288492 107778
rect 288440 107714 288492 107720
rect 288452 2938 288480 107714
rect 288820 106842 288848 110078
rect 289188 107794 289216 110078
rect 288544 106814 288848 106842
rect 288912 107766 289216 107794
rect 288544 4078 288572 106814
rect 288912 103514 288940 107766
rect 289924 107710 289952 110092
rect 290384 108594 290412 110092
rect 290372 108588 290424 108594
rect 290372 108530 290424 108536
rect 290752 107846 290780 110092
rect 290740 107840 290792 107846
rect 290740 107782 290792 107788
rect 291120 107778 291148 110092
rect 291304 110078 291594 110106
rect 291672 110078 291962 110106
rect 291108 107772 291160 107778
rect 291108 107714 291160 107720
rect 289084 107704 289136 107710
rect 289084 107646 289136 107652
rect 289912 107704 289964 107710
rect 289912 107646 289964 107652
rect 288636 103486 288940 103514
rect 288532 4072 288584 4078
rect 288532 4014 288584 4020
rect 288636 3058 288664 103486
rect 289096 4146 289124 107646
rect 291200 106820 291252 106826
rect 291200 106762 291252 106768
rect 289084 4140 289136 4146
rect 289084 4082 289136 4088
rect 290188 3596 290240 3602
rect 290188 3538 290240 3544
rect 288624 3052 288676 3058
rect 288624 2994 288676 3000
rect 288452 2910 289032 2938
rect 289004 480 289032 2910
rect 290200 480 290228 3538
rect 291212 3482 291240 106762
rect 291304 3602 291332 110078
rect 291672 106826 291700 110078
rect 292408 107710 292436 110092
rect 292592 110078 292790 110106
rect 292868 110078 293250 110106
rect 293328 110078 293618 110106
rect 292396 107704 292448 107710
rect 292396 107646 292448 107652
rect 291660 106820 291712 106826
rect 291660 106762 291712 106768
rect 292592 3602 292620 110078
rect 292672 107704 292724 107710
rect 292672 107646 292724 107652
rect 291292 3596 291344 3602
rect 291292 3538 291344 3544
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292684 3482 292712 107646
rect 292868 106842 292896 110078
rect 291212 3454 291424 3482
rect 291396 480 291424 3454
rect 292592 3454 292712 3482
rect 292776 106814 292896 106842
rect 292592 480 292620 3454
rect 292776 3058 292804 106814
rect 293328 103514 293356 110078
rect 292868 103486 293356 103514
rect 292868 3194 292896 103486
rect 293972 3738 294000 110092
rect 294064 110078 294446 110106
rect 293960 3732 294012 3738
rect 293960 3674 294012 3680
rect 293316 3596 293368 3602
rect 293316 3538 293368 3544
rect 292856 3188 292908 3194
rect 292856 3130 292908 3136
rect 292764 3052 292816 3058
rect 292764 2994 292816 3000
rect 287766 354 287878 480
rect 287440 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293328 354 293356 3538
rect 294064 3534 294092 110078
rect 294800 107710 294828 110092
rect 295260 108050 295288 110092
rect 295352 110078 295642 110106
rect 295720 110078 296010 110106
rect 296088 110078 296470 110106
rect 296838 110078 296944 110106
rect 295248 108044 295300 108050
rect 295248 107986 295300 107992
rect 294788 107704 294840 107710
rect 294788 107646 294840 107652
rect 295352 3942 295380 110078
rect 295432 106820 295484 106826
rect 295432 106762 295484 106768
rect 295340 3936 295392 3942
rect 295340 3878 295392 3884
rect 295444 3602 295472 106762
rect 295720 103514 295748 110078
rect 295984 107704 296036 107710
rect 295984 107646 296036 107652
rect 295536 103486 295748 103514
rect 295536 8974 295564 103486
rect 295524 8968 295576 8974
rect 295524 8910 295576 8916
rect 295996 4010 296024 107646
rect 296088 106826 296116 110078
rect 296720 108180 296772 108186
rect 296720 108122 296772 108128
rect 296076 106820 296128 106826
rect 296076 106762 296128 106768
rect 295984 4004 296036 4010
rect 295984 3946 296036 3952
rect 296732 3670 296760 108122
rect 296812 106820 296864 106826
rect 296812 106762 296864 106768
rect 296824 3806 296852 106762
rect 296812 3800 296864 3806
rect 296812 3742 296864 3748
rect 296720 3664 296772 3670
rect 296720 3606 296772 3612
rect 295432 3596 295484 3602
rect 295432 3538 295484 3544
rect 294052 3528 294104 3534
rect 294052 3470 294104 3476
rect 296916 3398 296944 110078
rect 297284 107710 297312 110092
rect 297376 110078 297666 110106
rect 297744 110078 298034 110106
rect 297376 108186 297404 110078
rect 297364 108180 297416 108186
rect 297364 108122 297416 108128
rect 297364 108044 297416 108050
rect 297364 107986 297416 107992
rect 297272 107704 297324 107710
rect 297272 107646 297324 107652
rect 297272 3732 297324 3738
rect 297272 3674 297324 3680
rect 296904 3392 296956 3398
rect 296904 3334 296956 3340
rect 296076 3188 296128 3194
rect 296076 3130 296128 3136
rect 294880 3052 294932 3058
rect 294880 2994 294932 3000
rect 294892 480 294920 2994
rect 296088 480 296116 3130
rect 297284 480 297312 3674
rect 297376 3262 297404 107986
rect 297744 106826 297772 110078
rect 298480 107778 298508 110092
rect 298572 110078 298862 110106
rect 299032 110078 299322 110106
rect 299584 110078 299690 110106
rect 298468 107772 298520 107778
rect 298468 107714 298520 107720
rect 297732 106820 297784 106826
rect 297732 106762 297784 106768
rect 298100 106820 298152 106826
rect 298100 106762 298152 106768
rect 298112 3670 298140 106762
rect 298572 103514 298600 110078
rect 299032 106826 299060 110078
rect 299020 106820 299072 106826
rect 299020 106762 299072 106768
rect 299480 103964 299532 103970
rect 299480 103906 299532 103912
rect 298204 103486 298600 103514
rect 298204 22778 298232 103486
rect 298192 22772 298244 22778
rect 298192 22714 298244 22720
rect 298100 3664 298152 3670
rect 298100 3606 298152 3612
rect 299492 3534 299520 103906
rect 299584 7750 299612 110078
rect 300044 108390 300072 110092
rect 300136 110078 300518 110106
rect 300886 110078 300992 110106
rect 300032 108384 300084 108390
rect 300032 108326 300084 108332
rect 300032 107704 300084 107710
rect 300032 107646 300084 107652
rect 300044 103514 300072 107646
rect 300136 103970 300164 110078
rect 300860 106888 300912 106894
rect 300860 106830 300912 106836
rect 300124 103964 300176 103970
rect 300124 103906 300176 103912
rect 300044 103486 300164 103514
rect 299572 7744 299624 7750
rect 299572 7686 299624 7692
rect 300136 4554 300164 103486
rect 300124 4548 300176 4554
rect 300124 4490 300176 4496
rect 299664 4004 299716 4010
rect 299664 3946 299716 3952
rect 298468 3528 298520 3534
rect 298468 3470 298520 3476
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 297364 3256 297416 3262
rect 297364 3198 297416 3204
rect 298480 480 298508 3470
rect 299676 480 299704 3946
rect 300872 3466 300900 106830
rect 300964 6254 300992 110078
rect 301148 110078 301346 110106
rect 301424 110078 301714 110106
rect 301792 110078 302174 110106
rect 302344 110078 302542 110106
rect 301044 106820 301096 106826
rect 301044 106762 301096 106768
rect 301056 11830 301084 106762
rect 301148 17270 301176 110078
rect 301424 106894 301452 110078
rect 301412 106888 301464 106894
rect 301412 106830 301464 106836
rect 301792 106826 301820 110078
rect 301780 106820 301832 106826
rect 301780 106762 301832 106768
rect 302240 106820 302292 106826
rect 302240 106762 302292 106768
rect 301136 17264 301188 17270
rect 301136 17206 301188 17212
rect 301044 11824 301096 11830
rect 301044 11766 301096 11772
rect 302252 10402 302280 106762
rect 302344 21622 302372 110078
rect 302896 108458 302924 110092
rect 303080 110078 303370 110106
rect 303632 110078 303738 110106
rect 303816 110078 304198 110106
rect 304276 110078 304566 110106
rect 302884 108452 302936 108458
rect 302884 108394 302936 108400
rect 302884 107772 302936 107778
rect 302884 107714 302936 107720
rect 302332 21616 302384 21622
rect 302332 21558 302384 21564
rect 302240 10396 302292 10402
rect 302240 10338 302292 10344
rect 302896 9042 302924 107714
rect 303080 106826 303108 110078
rect 303068 106820 303120 106826
rect 303068 106762 303120 106768
rect 302884 9036 302936 9042
rect 302884 8978 302936 8984
rect 303160 8968 303212 8974
rect 303160 8910 303212 8916
rect 300952 6248 301004 6254
rect 300952 6190 301004 6196
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 300860 3460 300912 3466
rect 300860 3402 300912 3408
rect 300768 3256 300820 3262
rect 300768 3198 300820 3204
rect 300780 480 300808 3198
rect 301976 480 302004 3878
rect 303172 480 303200 8910
rect 303632 6186 303660 110078
rect 303712 106820 303764 106826
rect 303712 106762 303764 106768
rect 303724 13190 303752 106762
rect 303816 15978 303844 110078
rect 304276 106826 304304 110078
rect 304920 108322 304948 110092
rect 305196 110078 305394 110106
rect 305472 110078 305762 110106
rect 305840 110078 306222 110106
rect 306484 110078 306590 110106
rect 306668 110078 306958 110106
rect 307128 110078 307418 110106
rect 304908 108316 304960 108322
rect 304908 108258 304960 108264
rect 305092 106888 305144 106894
rect 305092 106830 305144 106836
rect 304264 106820 304316 106826
rect 304264 106762 304316 106768
rect 305000 106820 305052 106826
rect 305000 106762 305052 106768
rect 303804 15972 303856 15978
rect 303804 15914 303856 15920
rect 303712 13184 303764 13190
rect 303712 13126 303764 13132
rect 305012 7682 305040 106762
rect 305104 10334 305132 106830
rect 305196 26926 305224 110078
rect 305472 106826 305500 110078
rect 305840 106894 305868 110078
rect 305828 106888 305880 106894
rect 305828 106830 305880 106836
rect 305460 106820 305512 106826
rect 305460 106762 305512 106768
rect 306380 106820 306432 106826
rect 306380 106762 306432 106768
rect 305184 26920 305236 26926
rect 305184 26862 305236 26868
rect 305092 10328 305144 10334
rect 305092 10270 305144 10276
rect 305000 7676 305052 7682
rect 305000 7618 305052 7624
rect 303620 6180 303672 6186
rect 303620 6122 303672 6128
rect 306392 4962 306420 106762
rect 306484 14618 306512 110078
rect 306668 103514 306696 110078
rect 307128 106826 307156 110078
rect 307116 106820 307168 106826
rect 307116 106762 307168 106768
rect 306576 103486 306696 103514
rect 306472 14612 306524 14618
rect 306472 14554 306524 14560
rect 306576 14482 306604 103486
rect 307772 31074 307800 110092
rect 308232 107710 308260 110092
rect 308600 107778 308628 110092
rect 308784 110078 309074 110106
rect 308588 107772 308640 107778
rect 308588 107714 308640 107720
rect 308220 107704 308272 107710
rect 308220 107646 308272 107652
rect 308784 103514 308812 110078
rect 309428 106962 309456 110092
rect 309520 110078 309810 110106
rect 309888 110078 310270 110106
rect 309416 106956 309468 106962
rect 309416 106898 309468 106904
rect 309520 106842 309548 110078
rect 309888 108474 309916 110078
rect 307864 103486 308812 103514
rect 309152 106814 309548 106842
rect 309612 108446 309916 108474
rect 307864 91798 307892 103486
rect 307852 91792 307904 91798
rect 307852 91734 307904 91740
rect 307760 31068 307812 31074
rect 307760 31010 307812 31016
rect 306564 14476 306616 14482
rect 306564 14418 306616 14424
rect 309152 6390 309180 106814
rect 309612 103514 309640 108446
rect 310624 108390 310652 110092
rect 310716 110078 311098 110106
rect 311176 110078 311466 110106
rect 311544 110078 311834 110106
rect 311912 110078 312294 110106
rect 312372 110078 312662 110106
rect 309784 108384 309836 108390
rect 309784 108326 309836 108332
rect 310612 108384 310664 108390
rect 310612 108326 310664 108332
rect 309244 103486 309640 103514
rect 309244 76566 309272 103486
rect 309232 76560 309284 76566
rect 309232 76502 309284 76508
rect 309796 9654 309824 108326
rect 309968 107704 310020 107710
rect 309968 107646 310020 107652
rect 309980 103514 310008 107646
rect 310716 106842 310744 110078
rect 310520 106820 310572 106826
rect 310520 106762 310572 106768
rect 310624 106814 310744 106842
rect 309888 103486 310008 103514
rect 309888 18698 309916 103486
rect 309876 18692 309928 18698
rect 309876 18634 309928 18640
rect 310532 11762 310560 106762
rect 310624 28490 310652 106814
rect 311176 106706 311204 110078
rect 311256 107772 311308 107778
rect 311256 107714 311308 107720
rect 310716 106678 311204 106706
rect 310716 61402 310744 106678
rect 311268 103514 311296 107714
rect 311544 106826 311572 110078
rect 311532 106820 311584 106826
rect 311532 106762 311584 106768
rect 311176 103486 311296 103514
rect 310704 61396 310756 61402
rect 310704 61338 310756 61344
rect 310612 28484 310664 28490
rect 310612 28426 310664 28432
rect 311176 25634 311204 103486
rect 311912 29646 311940 110078
rect 312372 99374 312400 110078
rect 313108 108594 313136 110092
rect 313292 110078 313490 110106
rect 313568 110078 313858 110106
rect 313936 110078 314318 110106
rect 313096 108588 313148 108594
rect 313096 108530 313148 108536
rect 312004 99346 312400 99374
rect 312004 73846 312032 99346
rect 311992 73840 312044 73846
rect 311992 73782 312044 73788
rect 311900 29640 311952 29646
rect 311900 29582 311952 29588
rect 311164 25628 311216 25634
rect 311164 25570 311216 25576
rect 310612 22772 310664 22778
rect 310612 22714 310664 22720
rect 310624 16574 310652 22714
rect 310624 16546 311480 16574
rect 310520 11756 310572 11762
rect 310520 11698 310572 11704
rect 309784 9648 309836 9654
rect 309784 9590 309836 9596
rect 310244 8968 310296 8974
rect 310244 8910 310296 8916
rect 309140 6384 309192 6390
rect 309140 6326 309192 6332
rect 306380 4956 306432 4962
rect 306380 4898 306432 4904
rect 306748 4548 306800 4554
rect 306748 4490 306800 4496
rect 304356 3596 304408 3602
rect 304356 3538 304408 3544
rect 304368 480 304396 3538
rect 305552 3392 305604 3398
rect 305552 3334 305604 3340
rect 305564 480 305592 3334
rect 306760 480 306788 4490
rect 309048 3800 309100 3806
rect 309048 3742 309100 3748
rect 307944 3664 307996 3670
rect 307944 3606 307996 3612
rect 307956 480 307984 3606
rect 309060 480 309088 3742
rect 310256 480 310284 8910
rect 311452 480 311480 16546
rect 313292 7614 313320 110078
rect 313372 104236 313424 104242
rect 313372 104178 313424 104184
rect 313384 15910 313412 104178
rect 313568 99374 313596 110078
rect 313936 104242 313964 110078
rect 314672 108866 314700 110092
rect 314764 110078 315146 110106
rect 315224 110078 315514 110106
rect 315592 110078 315882 110106
rect 316052 110078 316342 110106
rect 314660 108860 314712 108866
rect 314660 108802 314712 108808
rect 313924 104236 313976 104242
rect 313924 104178 313976 104184
rect 314660 104236 314712 104242
rect 314660 104178 314712 104184
rect 313476 99346 313596 99374
rect 313476 35222 313504 99346
rect 313464 35216 313516 35222
rect 313464 35158 313516 35164
rect 314672 22846 314700 104178
rect 314764 36582 314792 110078
rect 314844 108860 314896 108866
rect 314844 108802 314896 108808
rect 314856 66910 314884 108802
rect 315224 104242 315252 110078
rect 315304 108452 315356 108458
rect 315304 108394 315356 108400
rect 315212 104236 315264 104242
rect 315212 104178 315264 104184
rect 314844 66904 314896 66910
rect 314844 66846 314896 66852
rect 314752 36576 314804 36582
rect 314752 36518 314804 36524
rect 314660 22840 314712 22846
rect 314660 22782 314712 22788
rect 315316 17338 315344 108394
rect 315592 101454 315620 110078
rect 315580 101448 315632 101454
rect 315580 101390 315632 101396
rect 316052 37942 316080 110078
rect 316696 107710 316724 110092
rect 316788 110078 317170 110106
rect 317538 110078 317644 110106
rect 316684 107704 316736 107710
rect 316684 107646 316736 107652
rect 316788 99374 316816 110078
rect 317616 106274 317644 110078
rect 317432 106246 317644 106274
rect 317708 110078 317998 110106
rect 318076 110078 318366 110106
rect 318444 110078 318734 110106
rect 318812 110078 319194 110106
rect 319272 110078 319562 110106
rect 317432 104378 317460 106246
rect 317708 104514 317736 110078
rect 317512 104508 317564 104514
rect 317512 104450 317564 104456
rect 317696 104508 317748 104514
rect 317696 104450 317748 104456
rect 317420 104372 317472 104378
rect 317420 104314 317472 104320
rect 317420 104236 317472 104242
rect 317420 104178 317472 104184
rect 316144 99346 316816 99374
rect 316144 90370 316172 99346
rect 316132 90364 316184 90370
rect 316132 90306 316184 90312
rect 316040 37936 316092 37942
rect 316040 37878 316092 37884
rect 315304 17332 315356 17338
rect 315304 17274 315356 17280
rect 313372 15904 313424 15910
rect 313372 15846 313424 15852
rect 315028 9648 315080 9654
rect 315028 9590 315080 9596
rect 313832 7744 313884 7750
rect 313832 7686 313884 7692
rect 313280 7608 313332 7614
rect 313280 7550 313332 7556
rect 312636 3596 312688 3602
rect 312636 3538 312688 3544
rect 312648 480 312676 3538
rect 313844 480 313872 7686
rect 315040 480 315068 9590
rect 317432 9110 317460 104178
rect 317524 13122 317552 104450
rect 317604 104372 317656 104378
rect 317604 104314 317656 104320
rect 317616 50386 317644 104314
rect 318076 104242 318104 110078
rect 318064 104236 318116 104242
rect 318064 104178 318116 104184
rect 318444 99374 318472 110078
rect 317708 99346 318472 99374
rect 317708 58682 317736 99346
rect 317696 58676 317748 58682
rect 317696 58618 317748 58624
rect 317604 50380 317656 50386
rect 317604 50322 317656 50328
rect 317604 17264 317656 17270
rect 317604 17206 317656 17212
rect 317616 16574 317644 17206
rect 317616 16546 318104 16574
rect 317512 13116 317564 13122
rect 317512 13058 317564 13064
rect 317420 9104 317472 9110
rect 317420 9046 317472 9052
rect 317328 6248 317380 6254
rect 317328 6190 317380 6196
rect 316224 3528 316276 3534
rect 316224 3470 316276 3476
rect 316236 480 316264 3470
rect 317340 480 317368 6190
rect 293654 354 293766 480
rect 293328 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 318812 4894 318840 110078
rect 319272 99374 319300 110078
rect 320008 107982 320036 110092
rect 320192 110078 320390 110106
rect 320468 110078 320758 110106
rect 320836 110078 321218 110106
rect 319996 107976 320048 107982
rect 319996 107918 320048 107924
rect 319444 107704 319496 107710
rect 319444 107646 319496 107652
rect 318904 99346 319300 99374
rect 318904 9042 318932 99346
rect 319456 20058 319484 107646
rect 319444 20052 319496 20058
rect 319444 19994 319496 20000
rect 318892 9036 318944 9042
rect 318892 8978 318944 8984
rect 318800 4888 318852 4894
rect 318800 4830 318852 4836
rect 320192 4826 320220 110078
rect 320468 109034 320496 110078
rect 320284 109006 320496 109034
rect 320284 8974 320312 109006
rect 320836 99374 320864 110078
rect 321572 107710 321600 110092
rect 321664 110078 322046 110106
rect 322124 110078 322414 110106
rect 322492 110078 322782 110106
rect 322952 110078 323242 110106
rect 323320 110078 323610 110106
rect 323688 110078 324070 110106
rect 324438 110078 324544 110106
rect 321560 107704 321612 107710
rect 321560 107646 321612 107652
rect 321664 106978 321692 110078
rect 320376 99346 320864 99374
rect 321572 106950 321692 106978
rect 320376 51746 320404 99346
rect 320364 51740 320416 51746
rect 320364 51682 320416 51688
rect 321572 21486 321600 106950
rect 322124 106842 322152 110078
rect 321664 106814 322152 106842
rect 321664 53106 321692 106814
rect 322492 103514 322520 110078
rect 321756 103486 322520 103514
rect 321756 94518 321784 103486
rect 321744 94512 321796 94518
rect 321744 94454 321796 94460
rect 321652 53100 321704 53106
rect 321652 53042 321704 53048
rect 321652 21616 321704 21622
rect 321652 21558 321704 21564
rect 321560 21480 321612 21486
rect 321560 21422 321612 21428
rect 321664 16574 321692 21558
rect 321664 16546 322152 16574
rect 320456 11824 320508 11830
rect 320456 11766 320508 11772
rect 320272 8968 320324 8974
rect 320272 8910 320324 8916
rect 320180 4820 320232 4826
rect 320180 4762 320232 4768
rect 319720 3460 319772 3466
rect 319720 3402 319772 3408
rect 319732 480 319760 3402
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 11766
rect 322124 480 322152 16546
rect 322952 9450 322980 110078
rect 323032 105868 323084 105874
rect 323032 105810 323084 105816
rect 323044 24206 323072 105810
rect 323320 103514 323348 110078
rect 323584 107704 323636 107710
rect 323584 107646 323636 107652
rect 323136 103486 323348 103514
rect 323136 72486 323164 103486
rect 323124 72480 323176 72486
rect 323124 72422 323176 72428
rect 323032 24200 323084 24206
rect 323032 24142 323084 24148
rect 323596 17338 323624 107646
rect 323688 105874 323716 110078
rect 324320 106820 324372 106826
rect 324320 106762 324372 106768
rect 323676 105868 323728 105874
rect 323676 105810 323728 105816
rect 324332 32434 324360 106762
rect 324412 105596 324464 105602
rect 324412 105538 324464 105544
rect 324424 54602 324452 105538
rect 324516 55894 324544 110078
rect 324608 110078 324806 110106
rect 324884 110078 325266 110106
rect 325344 110078 325634 110106
rect 325712 110078 326094 110106
rect 324608 105602 324636 110078
rect 324596 105596 324648 105602
rect 324596 105538 324648 105544
rect 324884 103514 324912 110078
rect 325344 106826 325372 110078
rect 325332 106820 325384 106826
rect 325332 106762 325384 106768
rect 324608 103486 324912 103514
rect 324608 89010 324636 103486
rect 324596 89004 324648 89010
rect 324596 88946 324648 88952
rect 324504 55888 324556 55894
rect 324504 55830 324556 55836
rect 324412 54596 324464 54602
rect 324412 54538 324464 54544
rect 324320 32428 324372 32434
rect 324320 32370 324372 32376
rect 325712 25566 325740 110078
rect 326448 107710 326476 110092
rect 326540 110078 326922 110106
rect 327092 110078 327290 110106
rect 327368 110078 327658 110106
rect 327736 110078 328118 110106
rect 328486 110078 328684 110106
rect 326436 107704 326488 107710
rect 326436 107646 326488 107652
rect 326540 103514 326568 110078
rect 325804 103486 326568 103514
rect 325804 93294 325832 103486
rect 325792 93288 325844 93294
rect 325792 93230 325844 93236
rect 325700 25560 325752 25566
rect 325700 25502 325752 25508
rect 327092 22778 327120 110078
rect 327172 106820 327224 106826
rect 327172 106762 327224 106768
rect 327184 86290 327212 106762
rect 327368 103514 327396 110078
rect 327632 107976 327684 107982
rect 327632 107918 327684 107924
rect 327276 103486 327396 103514
rect 327644 103514 327672 107918
rect 327736 106826 327764 110078
rect 328460 108316 328512 108322
rect 328460 108258 328512 108264
rect 327816 107704 327868 107710
rect 327816 107646 327868 107652
rect 327724 106820 327776 106826
rect 327724 106762 327776 106768
rect 327644 103486 327764 103514
rect 327276 100094 327304 103486
rect 327264 100088 327316 100094
rect 327264 100030 327316 100036
rect 327172 86284 327224 86290
rect 327172 86226 327224 86232
rect 327080 22772 327132 22778
rect 327080 22714 327132 22720
rect 323032 17332 323084 17338
rect 323032 17274 323084 17280
rect 323584 17332 323636 17338
rect 323584 17274 323636 17280
rect 322940 9444 322992 9450
rect 322940 9386 322992 9392
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323044 354 323072 17274
rect 326344 15972 326396 15978
rect 326344 15914 326396 15920
rect 324412 10396 324464 10402
rect 324412 10338 324464 10344
rect 324424 480 324452 10338
rect 325608 6180 325660 6186
rect 325608 6122 325660 6128
rect 325620 480 325648 6122
rect 323278 354 323390 480
rect 323044 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 15914
rect 327736 14550 327764 103486
rect 327828 18630 327856 107646
rect 327816 18624 327868 18630
rect 327816 18566 327868 18572
rect 328472 16574 328500 108258
rect 328552 106820 328604 106826
rect 328552 106762 328604 106768
rect 328564 57322 328592 106762
rect 328656 60042 328684 110078
rect 328932 105738 328960 110092
rect 329024 110078 329314 110106
rect 329392 110078 329682 110106
rect 328920 105732 328972 105738
rect 328920 105674 328972 105680
rect 329024 103514 329052 110078
rect 329392 106826 329420 110078
rect 330128 108118 330156 110092
rect 330220 110078 330510 110106
rect 330680 110078 330970 110106
rect 330116 108112 330168 108118
rect 330116 108054 330168 108060
rect 329380 106820 329432 106826
rect 329380 106762 329432 106768
rect 329840 106820 329892 106826
rect 329840 106762 329892 106768
rect 328748 103486 329052 103514
rect 328748 96082 328776 103486
rect 328736 96076 328788 96082
rect 328736 96018 328788 96024
rect 329852 89078 329880 106762
rect 330220 103514 330248 110078
rect 330680 106826 330708 110078
rect 330668 106820 330720 106826
rect 330668 106762 330720 106768
rect 331220 106140 331272 106146
rect 331220 106082 331272 106088
rect 329944 103486 330248 103514
rect 329944 98802 329972 103486
rect 329932 98796 329984 98802
rect 329932 98738 329984 98744
rect 329840 89072 329892 89078
rect 329840 89014 329892 89020
rect 328644 60036 328696 60042
rect 328644 59978 328696 59984
rect 328552 57316 328604 57322
rect 328552 57258 328604 57264
rect 329840 26920 329892 26926
rect 329840 26862 329892 26868
rect 329852 16574 329880 26862
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 327724 14544 327776 14550
rect 327724 14486 327776 14492
rect 328000 13184 328052 13190
rect 328000 13126 328052 13132
rect 328012 480 328040 13126
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 331232 10878 331260 106082
rect 331324 104310 331352 110092
rect 331416 110078 331706 110106
rect 331784 110078 332166 110106
rect 332244 110078 332534 110106
rect 332704 110078 332994 110106
rect 331416 106146 331444 110078
rect 331404 106140 331456 106146
rect 331404 106082 331456 106088
rect 331312 104304 331364 104310
rect 331312 104246 331364 104252
rect 331784 104122 331812 110078
rect 331324 104094 331812 104122
rect 331324 62898 331352 104094
rect 332244 103514 332272 110078
rect 332600 106820 332652 106826
rect 332600 106762 332652 106768
rect 331416 103486 332272 103514
rect 331416 83570 331444 103486
rect 331404 83564 331456 83570
rect 331404 83506 331456 83512
rect 331312 62892 331364 62898
rect 331312 62834 331364 62840
rect 331220 10872 331272 10878
rect 331220 10814 331272 10820
rect 331588 7676 331640 7682
rect 331588 7618 331640 7624
rect 331600 480 331628 7618
rect 332612 6322 332640 106762
rect 332704 10810 332732 110078
rect 333348 108458 333376 110092
rect 333440 110078 333730 110106
rect 333992 110078 334190 110106
rect 334268 110078 334558 110106
rect 334636 110078 335018 110106
rect 335386 110078 335492 110106
rect 333336 108452 333388 108458
rect 333336 108394 333388 108400
rect 333244 108384 333296 108390
rect 333244 108326 333296 108332
rect 332692 10804 332744 10810
rect 332692 10746 332744 10752
rect 332692 10328 332744 10334
rect 332692 10270 332744 10276
rect 332600 6316 332652 6322
rect 332600 6258 332652 6264
rect 332704 480 332732 10270
rect 333256 7682 333284 108326
rect 333440 106826 333468 110078
rect 333428 106820 333480 106826
rect 333428 106762 333480 106768
rect 333888 14612 333940 14618
rect 333888 14554 333940 14560
rect 333244 7676 333296 7682
rect 333244 7618 333296 7624
rect 333900 480 333928 14554
rect 333992 10742 334020 110078
rect 334268 106842 334296 110078
rect 334084 106814 334296 106842
rect 334084 19990 334112 106814
rect 334636 103514 334664 110078
rect 335360 106888 335412 106894
rect 335360 106830 335412 106836
rect 334176 103486 334664 103514
rect 334176 82210 334204 103486
rect 334164 82204 334216 82210
rect 334164 82146 334216 82152
rect 334072 19984 334124 19990
rect 334072 19926 334124 19932
rect 334624 14476 334676 14482
rect 334624 14418 334676 14424
rect 333980 10736 334032 10742
rect 333980 10678 334032 10684
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 14418
rect 335372 6254 335400 106830
rect 335464 10674 335492 110078
rect 335648 110078 335846 110106
rect 335924 110078 336214 110106
rect 336292 110078 336582 110106
rect 336936 110078 337042 110106
rect 337120 110078 337410 110106
rect 337488 110078 337870 110106
rect 338132 110078 338238 110106
rect 338316 110078 338606 110106
rect 338776 110078 339066 110106
rect 335544 106820 335596 106826
rect 335544 106762 335596 106768
rect 335452 10668 335504 10674
rect 335452 10610 335504 10616
rect 335556 10606 335584 106762
rect 335648 93226 335676 110078
rect 335924 106894 335952 110078
rect 335912 106888 335964 106894
rect 335912 106830 335964 106836
rect 336292 106826 336320 110078
rect 336280 106820 336332 106826
rect 336280 106762 336332 106768
rect 336740 106820 336792 106826
rect 336740 106762 336792 106768
rect 335636 93220 335688 93226
rect 335636 93162 335688 93168
rect 335544 10600 335596 10606
rect 335544 10542 335596 10548
rect 335360 6248 335412 6254
rect 335360 6190 335412 6196
rect 336752 6186 336780 106762
rect 336832 106684 336884 106690
rect 336832 106626 336884 106632
rect 336844 10538 336872 106626
rect 336936 96014 336964 110078
rect 337120 106826 337148 110078
rect 337384 108112 337436 108118
rect 337384 108054 337436 108060
rect 337108 106820 337160 106826
rect 337108 106762 337160 106768
rect 336924 96008 336976 96014
rect 336924 95950 336976 95956
rect 337396 84930 337424 108054
rect 337488 106690 337516 110078
rect 337476 106684 337528 106690
rect 337476 106626 337528 106632
rect 337384 84924 337436 84930
rect 337384 84866 337436 84872
rect 336924 31068 336976 31074
rect 336924 31010 336976 31016
rect 336936 16574 336964 31010
rect 336936 16546 337056 16574
rect 336832 10532 336884 10538
rect 336832 10474 336884 10480
rect 336740 6180 336792 6186
rect 336740 6122 336792 6128
rect 336280 4956 336332 4962
rect 336280 4898 336332 4904
rect 336292 480 336320 4898
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338132 3262 338160 110078
rect 338212 106820 338264 106826
rect 338212 106762 338264 106768
rect 338224 10470 338252 106762
rect 338316 80782 338344 110078
rect 338672 108452 338724 108458
rect 338672 108394 338724 108400
rect 338684 103514 338712 108394
rect 338776 106826 338804 110078
rect 339420 108662 339448 110092
rect 339408 108656 339460 108662
rect 339408 108598 339460 108604
rect 339880 107098 339908 110092
rect 339972 110078 340262 110106
rect 340340 110078 340630 110106
rect 339868 107092 339920 107098
rect 339868 107034 339920 107040
rect 338764 106820 338816 106826
rect 338764 106762 338816 106768
rect 339500 106820 339552 106826
rect 339500 106762 339552 106768
rect 338684 103486 338804 103514
rect 338304 80776 338356 80782
rect 338304 80718 338356 80724
rect 338776 29714 338804 103486
rect 338764 29708 338816 29714
rect 338764 29650 338816 29656
rect 338304 18692 338356 18698
rect 338304 18634 338356 18640
rect 338316 16574 338344 18634
rect 338316 16546 338712 16574
rect 338212 10464 338264 10470
rect 338212 10406 338264 10412
rect 338120 3256 338172 3262
rect 338120 3198 338172 3204
rect 338684 480 338712 16546
rect 339512 3330 339540 106762
rect 339972 103514 340000 110078
rect 340340 106826 340368 110078
rect 340880 106956 340932 106962
rect 340880 106898 340932 106904
rect 340328 106820 340380 106826
rect 340328 106762 340380 106768
rect 339604 103486 340000 103514
rect 339604 10402 339632 103486
rect 339684 25628 339736 25634
rect 339684 25570 339736 25576
rect 339592 10396 339644 10402
rect 339592 10338 339644 10344
rect 339500 3324 339552 3330
rect 339500 3266 339552 3272
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339696 354 339724 25570
rect 340892 3534 340920 106898
rect 340972 91792 341024 91798
rect 340972 91734 341024 91740
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 340984 480 341012 91734
rect 341076 26994 341104 110092
rect 341168 110078 341458 110106
rect 341168 91866 341196 110078
rect 341904 108458 341932 110092
rect 342286 110078 342484 110106
rect 341892 108452 341944 108458
rect 341892 108394 341944 108400
rect 342456 106978 342484 110078
rect 342640 110078 342746 110106
rect 342824 110078 343114 110106
rect 343192 110078 343482 110106
rect 343652 110078 343942 110106
rect 342456 106950 342576 106978
rect 342260 106888 342312 106894
rect 342260 106830 342312 106836
rect 341156 91860 341208 91866
rect 341156 91802 341208 91808
rect 341064 26988 341116 26994
rect 341064 26930 341116 26936
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 342272 3398 342300 106830
rect 342444 106820 342496 106826
rect 342444 106762 342496 106768
rect 342352 106752 342404 106758
rect 342352 106694 342404 106700
rect 342364 10334 342392 106694
rect 342456 78062 342484 106762
rect 342548 79422 342576 106950
rect 342640 106758 342668 110078
rect 342824 106894 342852 110078
rect 342812 106888 342864 106894
rect 342812 106830 342864 106836
rect 343192 106826 343220 110078
rect 343180 106820 343232 106826
rect 343180 106762 343232 106768
rect 342628 106752 342680 106758
rect 342628 106694 342680 106700
rect 343652 97374 343680 110078
rect 344296 108390 344324 110092
rect 344388 110078 344770 110106
rect 344284 108384 344336 108390
rect 344284 108326 344336 108332
rect 344388 103514 344416 110078
rect 343744 103486 344416 103514
rect 343640 97368 343692 97374
rect 343640 97310 343692 97316
rect 342536 79416 342588 79422
rect 342536 79358 342588 79364
rect 342444 78056 342496 78062
rect 342444 77998 342496 78004
rect 343744 76634 343772 103486
rect 343732 76628 343784 76634
rect 343732 76570 343784 76576
rect 343640 76560 343692 76566
rect 343640 76502 343692 76508
rect 343652 16574 343680 76502
rect 343652 16546 344600 16574
rect 342352 10328 342404 10334
rect 342352 10270 342404 10276
rect 343364 6384 343416 6390
rect 343364 6326 343416 6332
rect 342260 3392 342312 3398
rect 342260 3334 342312 3340
rect 343376 480 343404 6326
rect 344572 480 344600 16546
rect 345032 4146 345060 110162
rect 345138 110078 345336 110106
rect 345112 106888 345164 106894
rect 345112 106830 345164 106836
rect 345124 33862 345152 106830
rect 345204 106820 345256 106826
rect 345204 106762 345256 106768
rect 345216 75274 345244 106762
rect 345308 87718 345336 110078
rect 345584 110078 345966 110106
rect 346044 110078 346334 110106
rect 345584 106826 345612 110078
rect 346044 106894 346072 110078
rect 346780 108322 346808 110092
rect 346872 110078 347162 110106
rect 347240 110078 347530 110106
rect 347792 110078 347990 110106
rect 346768 108316 346820 108322
rect 346768 108258 346820 108264
rect 346032 106888 346084 106894
rect 346872 106842 346900 110078
rect 347240 108202 347268 110078
rect 346032 106830 346084 106836
rect 345572 106820 345624 106826
rect 345572 106762 345624 106768
rect 346412 106814 346900 106842
rect 346964 108174 347268 108202
rect 345296 87712 345348 87718
rect 345296 87654 345348 87660
rect 345204 75268 345256 75274
rect 345204 75210 345256 75216
rect 345112 33856 345164 33862
rect 345112 33798 345164 33804
rect 346412 28354 346440 106814
rect 346964 103514 346992 108174
rect 347044 108112 347096 108118
rect 347044 108054 347096 108060
rect 346504 103486 346992 103514
rect 346504 49094 346532 103486
rect 346492 49088 346544 49094
rect 346492 49030 346544 49036
rect 346492 28484 346544 28490
rect 346492 28426 346544 28432
rect 346400 28348 346452 28354
rect 346400 28290 346452 28296
rect 346504 16574 346532 28426
rect 346504 16546 346992 16574
rect 345756 7676 345808 7682
rect 345756 7618 345808 7624
rect 345020 4140 345072 4146
rect 345020 4082 345072 4088
rect 345768 480 345796 7618
rect 346964 480 346992 16546
rect 347056 4214 347084 108054
rect 347044 4208 347096 4214
rect 347044 4150 347096 4156
rect 347792 4078 347820 110078
rect 348344 107710 348372 110092
rect 348436 110078 348818 110106
rect 349186 110078 349292 110106
rect 348332 107704 348384 107710
rect 348332 107646 348384 107652
rect 348436 103514 348464 110078
rect 349160 106820 349212 106826
rect 349160 106762 349212 106768
rect 347884 103486 348464 103514
rect 347884 100026 347912 103486
rect 347872 100020 347924 100026
rect 347872 99962 347924 99968
rect 347872 61396 347924 61402
rect 347872 61338 347924 61344
rect 347884 16574 347912 61338
rect 347884 16546 348096 16574
rect 347780 4072 347832 4078
rect 347780 4014 347832 4020
rect 348068 480 348096 16546
rect 349172 3942 349200 106762
rect 349264 4010 349292 110078
rect 349344 106888 349396 106894
rect 349344 106830 349396 106836
rect 349356 47666 349384 106830
rect 349540 103578 349568 110092
rect 349632 110078 350014 110106
rect 350092 110078 350382 110106
rect 350644 110078 350842 110106
rect 350920 110078 351210 110106
rect 351288 110078 351670 110106
rect 349632 106894 349660 110078
rect 349620 106888 349672 106894
rect 349620 106830 349672 106836
rect 350092 106826 350120 110078
rect 350080 106820 350132 106826
rect 350080 106762 350132 106768
rect 350540 106820 350592 106826
rect 350540 106762 350592 106768
rect 349448 103550 349568 103578
rect 349448 102882 349476 103550
rect 349436 102876 349488 102882
rect 349436 102818 349488 102824
rect 349344 47660 349396 47666
rect 349344 47602 349396 47608
rect 349344 29640 349396 29646
rect 349344 29582 349396 29588
rect 349356 16574 349384 29582
rect 349356 16546 350488 16574
rect 349344 11756 349396 11762
rect 349344 11698 349396 11704
rect 349252 4004 349304 4010
rect 349252 3946 349304 3952
rect 349160 3936 349212 3942
rect 349160 3878 349212 3884
rect 349356 3482 349384 11698
rect 349264 3454 349384 3482
rect 349264 480 349292 3454
rect 350460 480 350488 16546
rect 350552 3874 350580 106762
rect 350644 7818 350672 110078
rect 350920 103514 350948 110078
rect 351184 107704 351236 107710
rect 351184 107646 351236 107652
rect 350736 103486 350948 103514
rect 350736 90438 350764 103486
rect 350724 90432 350776 90438
rect 350724 90374 350776 90380
rect 351196 73914 351224 107646
rect 351288 106826 351316 110078
rect 352024 107710 352052 110092
rect 352116 110078 352406 110106
rect 352576 110078 352866 110106
rect 352944 110078 353234 110106
rect 353496 110078 353694 110106
rect 353772 110078 354062 110106
rect 354140 110078 354430 110106
rect 352012 107704 352064 107710
rect 352012 107646 352064 107652
rect 351276 106820 351328 106826
rect 351276 106762 351328 106768
rect 352012 106820 352064 106826
rect 352012 106762 352064 106768
rect 351920 104780 351972 104786
rect 351920 104722 351972 104728
rect 351184 73908 351236 73914
rect 351184 73850 351236 73856
rect 350724 73840 350776 73846
rect 350724 73782 350776 73788
rect 350736 16574 350764 73782
rect 350736 16546 351224 16574
rect 350632 7812 350684 7818
rect 350632 7754 350684 7760
rect 350540 3868 350592 3874
rect 350540 3810 350592 3816
rect 339838 354 339950 480
rect 339696 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 351932 3806 351960 104722
rect 352024 69766 352052 106762
rect 352116 94586 352144 110078
rect 352576 104786 352604 110078
rect 352944 106826 352972 110078
rect 353392 106888 353444 106894
rect 353392 106830 353444 106836
rect 352932 106820 352984 106826
rect 352932 106762 352984 106768
rect 353300 106820 353352 106826
rect 353300 106762 353352 106768
rect 352564 104780 352616 104786
rect 352564 104722 352616 104728
rect 352104 94580 352156 94586
rect 352104 94522 352156 94528
rect 352012 69760 352064 69766
rect 352012 69702 352064 69708
rect 352840 4208 352892 4214
rect 352840 4150 352892 4156
rect 351920 3800 351972 3806
rect 351920 3742 351972 3748
rect 352852 480 352880 4150
rect 353312 3738 353340 106762
rect 353404 7750 353432 106830
rect 353496 46238 353524 110078
rect 353772 106826 353800 110078
rect 353944 107704 353996 107710
rect 353944 107646 353996 107652
rect 353760 106820 353812 106826
rect 353760 106762 353812 106768
rect 353956 71126 353984 107646
rect 354140 106894 354168 110078
rect 354128 106888 354180 106894
rect 354128 106830 354180 106836
rect 354772 106888 354824 106894
rect 354772 106830 354824 106836
rect 354680 106820 354732 106826
rect 354680 106762 354732 106768
rect 353944 71120 353996 71126
rect 353944 71062 353996 71068
rect 353484 46232 353536 46238
rect 353484 46174 353536 46180
rect 353392 7744 353444 7750
rect 353392 7686 353444 7692
rect 354036 7608 354088 7614
rect 354036 7550 354088 7556
rect 353300 3732 353352 3738
rect 353300 3674 353352 3680
rect 354048 480 354076 7550
rect 354692 3670 354720 106762
rect 354784 7682 354812 106830
rect 354876 11898 354904 110092
rect 354968 110078 355258 110106
rect 355336 110078 355718 110106
rect 356086 110078 356192 110106
rect 354968 106826 354996 110078
rect 355336 106894 355364 110078
rect 355324 106888 355376 106894
rect 355324 106830 355376 106836
rect 354956 106820 355008 106826
rect 354956 106762 355008 106768
rect 356060 106820 356112 106826
rect 356060 106762 356112 106768
rect 354956 35216 355008 35222
rect 354956 35158 355008 35164
rect 354968 16574 354996 35158
rect 354968 16546 355272 16574
rect 354864 11892 354916 11898
rect 354864 11834 354916 11840
rect 354772 7676 354824 7682
rect 354772 7618 354824 7624
rect 354680 3664 354732 3670
rect 354680 3606 354732 3612
rect 355244 480 355272 16546
rect 356072 3602 356100 106762
rect 356164 44878 356192 110078
rect 356256 110078 356454 110106
rect 356256 106826 356284 110078
rect 356900 107030 356928 110092
rect 356992 110078 357282 110106
rect 357544 110078 357742 110106
rect 356888 107024 356940 107030
rect 356888 106966 356940 106972
rect 356244 106820 356296 106826
rect 356244 106762 356296 106768
rect 356992 103514 357020 110078
rect 356256 103486 357020 103514
rect 356256 68406 356284 103486
rect 356244 68400 356296 68406
rect 356244 68342 356296 68348
rect 357440 66904 357492 66910
rect 357440 66846 357492 66852
rect 356152 44872 356204 44878
rect 356152 44814 356204 44820
rect 356336 15904 356388 15910
rect 356336 15846 356388 15852
rect 356060 3596 356112 3602
rect 356060 3538 356112 3544
rect 356348 480 356376 15846
rect 357452 3346 357480 66846
rect 357544 43450 357572 110078
rect 358096 105670 358124 110092
rect 358188 110078 358478 110106
rect 358084 105664 358136 105670
rect 358084 105606 358136 105612
rect 358188 103514 358216 110078
rect 358820 106820 358872 106826
rect 358820 106762 358872 106768
rect 357636 103486 358216 103514
rect 357636 66910 357664 103486
rect 357624 66904 357676 66910
rect 357624 66846 357676 66852
rect 357532 43444 357584 43450
rect 357532 43386 357584 43392
rect 357532 36576 357584 36582
rect 357532 36518 357584 36524
rect 357544 3534 357572 36518
rect 358832 35222 358860 106762
rect 358924 42090 358952 110092
rect 359292 104242 359320 110092
rect 359384 110078 359766 110106
rect 359844 110078 360134 110106
rect 360304 110078 360594 110106
rect 360672 110078 360962 110106
rect 361040 110078 361330 110106
rect 359280 104236 359332 104242
rect 359280 104178 359332 104184
rect 359384 103514 359412 110078
rect 359844 106826 359872 110078
rect 359832 106820 359884 106826
rect 359832 106762 359884 106768
rect 359016 103486 359412 103514
rect 359016 65550 359044 103486
rect 360304 102814 360332 110078
rect 360672 109034 360700 110078
rect 360396 109006 360700 109034
rect 360292 102808 360344 102814
rect 360292 102750 360344 102756
rect 360396 102626 360424 109006
rect 360212 102598 360424 102626
rect 359004 65544 359056 65550
rect 359004 65486 359056 65492
rect 358912 42084 358964 42090
rect 358912 42026 358964 42032
rect 358820 35216 358872 35222
rect 358820 35158 358872 35164
rect 358820 22840 358872 22846
rect 358820 22782 358872 22788
rect 358832 16574 358860 22782
rect 358832 16546 359504 16574
rect 357532 3528 357584 3534
rect 357532 3470 357584 3476
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 357452 3318 357572 3346
rect 357544 480 357572 3318
rect 358740 480 358768 3470
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 360212 7614 360240 102598
rect 360292 101448 360344 101454
rect 360292 101390 360344 101396
rect 360200 7608 360252 7614
rect 360200 7550 360252 7556
rect 360304 6914 360332 101390
rect 361040 99374 361068 110078
rect 361580 102196 361632 102202
rect 361580 102138 361632 102144
rect 360396 99346 361068 99374
rect 360396 11830 360424 99346
rect 361592 36582 361620 102138
rect 361776 101522 361804 110092
rect 361868 110078 362158 110106
rect 362328 110078 362618 110106
rect 362986 110078 363276 110106
rect 361764 101516 361816 101522
rect 361764 101458 361816 101464
rect 361868 99374 361896 110078
rect 362328 102202 362356 110078
rect 363248 105466 363276 110078
rect 363236 105460 363288 105466
rect 363236 105402 363288 105408
rect 363052 104168 363104 104174
rect 363052 104110 363104 104116
rect 362960 104100 363012 104106
rect 362960 104042 363012 104048
rect 362316 102196 362368 102202
rect 362316 102138 362368 102144
rect 361684 99346 361896 99374
rect 361684 84862 361712 99346
rect 361672 84856 361724 84862
rect 361672 84798 361724 84804
rect 361672 37936 361724 37942
rect 361672 37878 361724 37884
rect 361580 36576 361632 36582
rect 361580 36518 361632 36524
rect 361684 16574 361712 37878
rect 362972 17270 363000 104042
rect 363064 40730 363092 104110
rect 363340 96614 363368 110092
rect 363432 110078 363814 110106
rect 363892 110078 364182 110106
rect 363432 104174 363460 110078
rect 363512 105460 363564 105466
rect 363512 105402 363564 105408
rect 363420 104168 363472 104174
rect 363420 104110 363472 104116
rect 363524 98734 363552 105402
rect 363892 104106 363920 110078
rect 364340 104168 364392 104174
rect 364340 104110 364392 104116
rect 363880 104100 363932 104106
rect 363880 104042 363932 104048
rect 363512 98728 363564 98734
rect 363512 98670 363564 98676
rect 363156 96586 363368 96614
rect 363156 64190 363184 96586
rect 363144 64184 363196 64190
rect 363144 64126 363196 64132
rect 363052 40724 363104 40730
rect 363052 40666 363104 40672
rect 363052 20052 363104 20058
rect 363052 19994 363104 20000
rect 362960 17264 363012 17270
rect 362960 17206 363012 17212
rect 363064 16574 363092 19994
rect 361684 16546 361896 16574
rect 363064 16546 363552 16574
rect 360384 11824 360436 11830
rect 360384 11766 360436 11772
rect 360304 6886 361160 6914
rect 361132 480 361160 6886
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364352 11762 364380 104110
rect 364432 104100 364484 104106
rect 364432 104042 364484 104048
rect 364444 14482 364472 104042
rect 364524 90364 364576 90370
rect 364524 90306 364576 90312
rect 364536 16574 364564 90306
rect 364628 62830 364656 110092
rect 364720 110078 365010 110106
rect 365088 110078 365378 110106
rect 364720 104174 364748 110078
rect 364708 104168 364760 104174
rect 364708 104110 364760 104116
rect 365088 104106 365116 110078
rect 365824 107778 365852 110092
rect 365916 110078 366206 110106
rect 365812 107772 365864 107778
rect 365812 107714 365864 107720
rect 365916 104258 365944 110078
rect 366652 107710 366680 110092
rect 366744 110078 367034 110106
rect 367204 110078 367494 110106
rect 367572 110078 367862 110106
rect 367940 110078 368230 110106
rect 368584 110078 368690 110106
rect 368768 110078 369058 110106
rect 369136 110078 369518 110106
rect 369886 110078 369992 110106
rect 366640 107704 366692 107710
rect 366640 107646 366692 107652
rect 365732 104230 365944 104258
rect 365076 104100 365128 104106
rect 365076 104042 365128 104048
rect 364616 62824 364668 62830
rect 364616 62766 364668 62772
rect 365732 39370 365760 104230
rect 366744 99374 366772 110078
rect 367100 104168 367152 104174
rect 367100 104110 367152 104116
rect 365824 99346 366772 99374
rect 365824 82142 365852 99346
rect 365812 82136 365864 82142
rect 365812 82078 365864 82084
rect 365812 50380 365864 50386
rect 365812 50322 365864 50328
rect 365720 39364 365772 39370
rect 365720 39306 365772 39312
rect 364536 16546 364656 16574
rect 364432 14476 364484 14482
rect 364432 14418 364484 14424
rect 364340 11756 364392 11762
rect 364340 11698 364392 11704
rect 364628 480 364656 16546
rect 365720 13116 365772 13122
rect 365720 13058 365772 13064
rect 365732 3466 365760 13058
rect 365720 3460 365772 3466
rect 365720 3402 365772 3408
rect 365824 480 365852 50322
rect 367112 5166 367140 104110
rect 367204 13258 367232 110078
rect 367572 104174 367600 110078
rect 367940 109034 367968 110078
rect 367664 109006 367968 109034
rect 367560 104168 367612 104174
rect 367560 104110 367612 104116
rect 367664 99374 367692 109006
rect 367744 107704 367796 107710
rect 367744 107646 367796 107652
rect 367296 99346 367692 99374
rect 367296 61402 367324 99346
rect 367756 97306 367784 107646
rect 368584 106274 368612 110078
rect 368768 109034 368796 110078
rect 369136 109034 369164 110078
rect 368492 106246 368612 106274
rect 368676 109006 368796 109034
rect 369044 109006 369164 109034
rect 368492 101538 368520 106246
rect 368492 101510 368612 101538
rect 368480 101448 368532 101454
rect 368480 101390 368532 101396
rect 367744 97300 367796 97306
rect 367744 97242 367796 97248
rect 367284 61396 367336 61402
rect 367284 61338 367336 61344
rect 368492 15910 368520 101390
rect 368584 37942 368612 101510
rect 368676 101454 368704 109006
rect 368664 101448 368716 101454
rect 368664 101390 368716 101396
rect 369044 99374 369072 109006
rect 369124 107772 369176 107778
rect 369124 107714 369176 107720
rect 368768 99346 369072 99374
rect 368768 58682 368796 99346
rect 369136 83502 369164 107714
rect 369860 104168 369912 104174
rect 369860 104110 369912 104116
rect 369124 83496 369176 83502
rect 369124 83438 369176 83444
rect 369872 77994 369900 104110
rect 369964 79354 369992 110078
rect 370240 108594 370268 110092
rect 370332 110078 370714 110106
rect 370792 110078 371082 110106
rect 371344 110078 371542 110106
rect 371620 110078 371910 110106
rect 371988 110078 372278 110106
rect 370228 108588 370280 108594
rect 370228 108530 370280 108536
rect 370332 99374 370360 110078
rect 370792 104174 370820 110078
rect 370780 104168 370832 104174
rect 370780 104110 370832 104116
rect 371240 104168 371292 104174
rect 371240 104110 371292 104116
rect 370056 99346 370360 99374
rect 370056 80714 370084 99346
rect 370044 80708 370096 80714
rect 370044 80650 370096 80656
rect 369952 79348 370004 79354
rect 369952 79290 370004 79296
rect 369860 77988 369912 77994
rect 369860 77930 369912 77936
rect 368664 58676 368716 58682
rect 368664 58618 368716 58624
rect 368756 58676 368808 58682
rect 368756 58618 368808 58624
rect 368572 37936 368624 37942
rect 368572 37878 368624 37884
rect 368676 16574 368704 58618
rect 368676 16546 369440 16574
rect 368480 15904 368532 15910
rect 368480 15846 368532 15852
rect 367192 13252 367244 13258
rect 367192 13194 367244 13200
rect 368204 9104 368256 9110
rect 368204 9046 368256 9052
rect 367100 5160 367152 5166
rect 367100 5102 367152 5108
rect 367008 3460 367060 3466
rect 367008 3402 367060 3408
rect 367020 480 367048 3402
rect 368216 480 368244 9046
rect 369412 480 369440 16546
rect 371252 13190 371280 104110
rect 371344 21418 371372 110078
rect 371620 99374 371648 110078
rect 371988 104174 372016 110078
rect 371976 104168 372028 104174
rect 371976 104110 372028 104116
rect 372620 104168 372672 104174
rect 372620 104110 372672 104116
rect 371436 99346 371648 99374
rect 371436 31074 371464 99346
rect 371424 31068 371476 31074
rect 371424 31010 371476 31016
rect 371332 21412 371384 21418
rect 371332 21354 371384 21360
rect 371240 13184 371292 13190
rect 371240 13126 371292 13132
rect 371700 9036 371752 9042
rect 371700 8978 371752 8984
rect 370596 4888 370648 4894
rect 370596 4830 370648 4836
rect 370608 480 370636 4830
rect 371712 480 371740 8978
rect 372632 5030 372660 104110
rect 372724 5098 372752 110092
rect 372816 110078 373106 110106
rect 373184 110078 373566 110106
rect 373644 110078 373934 110106
rect 374104 110078 374302 110106
rect 374380 110078 374762 110106
rect 374840 110078 375130 110106
rect 375484 110078 375590 110106
rect 375668 110078 375958 110106
rect 376128 110078 376418 110106
rect 376786 110078 376892 110106
rect 372816 9382 372844 110078
rect 373184 99374 373212 110078
rect 373644 104174 373672 110078
rect 373632 104168 373684 104174
rect 373632 104110 373684 104116
rect 374000 104168 374052 104174
rect 374000 104110 374052 104116
rect 372908 99346 373212 99374
rect 372908 76566 372936 99346
rect 372896 76560 372948 76566
rect 372896 76502 372948 76508
rect 372896 14544 372948 14550
rect 372896 14486 372948 14492
rect 372804 9376 372856 9382
rect 372804 9318 372856 9324
rect 372712 5092 372764 5098
rect 372712 5034 372764 5040
rect 372620 5024 372672 5030
rect 372620 4966 372672 4972
rect 372908 480 372936 14486
rect 374012 4962 374040 104110
rect 374104 9314 374132 110078
rect 374380 99374 374408 110078
rect 374840 104174 374868 110078
rect 374828 104168 374880 104174
rect 374828 104110 374880 104116
rect 375484 101454 375512 110078
rect 375668 109034 375696 110078
rect 375576 109006 375696 109034
rect 375472 101448 375524 101454
rect 375472 101390 375524 101396
rect 375576 101266 375604 109006
rect 374196 99346 374408 99374
rect 375392 101238 375604 101266
rect 374196 13122 374224 99346
rect 375392 75206 375420 101238
rect 376128 99374 376156 110078
rect 376760 104168 376812 104174
rect 376760 104110 376812 104116
rect 375484 99346 376156 99374
rect 375484 95946 375512 99346
rect 375472 95940 375524 95946
rect 375472 95882 375524 95888
rect 375380 75200 375432 75206
rect 375380 75142 375432 75148
rect 375380 51740 375432 51746
rect 375380 51682 375432 51688
rect 375392 16574 375420 51682
rect 375392 16546 376064 16574
rect 374184 13116 374236 13122
rect 374184 13058 374236 13064
rect 374092 9308 374144 9314
rect 374092 9250 374144 9256
rect 375288 8968 375340 8974
rect 375288 8910 375340 8916
rect 374000 4956 374052 4962
rect 374000 4898 374052 4904
rect 374092 4820 374144 4826
rect 374092 4762 374144 4768
rect 374104 480 374132 4762
rect 375300 480 375328 8910
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 376772 4894 376800 104110
rect 376864 9246 376892 110078
rect 377140 104106 377168 110092
rect 377232 110078 377614 110106
rect 377692 110078 377982 110106
rect 378336 110078 378442 110106
rect 378520 110078 378810 110106
rect 378888 110078 379178 110106
rect 377232 104174 377260 110078
rect 377220 104168 377272 104174
rect 377220 104110 377272 104116
rect 377128 104100 377180 104106
rect 377128 104042 377180 104048
rect 377692 99374 377720 110078
rect 378336 106274 378364 110078
rect 378520 109034 378548 110078
rect 378244 106246 378364 106274
rect 378428 109006 378548 109034
rect 378140 104508 378192 104514
rect 378140 104450 378192 104456
rect 376956 99346 377720 99374
rect 376852 9240 376904 9246
rect 376852 9182 376904 9188
rect 376956 9178 376984 99346
rect 377036 17332 377088 17338
rect 377036 17274 377088 17280
rect 377048 16574 377076 17274
rect 377048 16546 377720 16574
rect 376944 9172 376996 9178
rect 376944 9114 376996 9120
rect 376760 4888 376812 4894
rect 376760 4830 376812 4836
rect 377692 480 377720 16546
rect 378152 4826 378180 104450
rect 378244 104258 378272 106246
rect 378428 104514 378456 109006
rect 378416 104508 378468 104514
rect 378416 104450 378468 104456
rect 378244 104230 378364 104258
rect 378232 104168 378284 104174
rect 378232 104110 378284 104116
rect 378244 9110 378272 104110
rect 378336 73846 378364 104230
rect 378888 104174 378916 110078
rect 379624 106962 379652 110092
rect 379992 107710 380020 110092
rect 379980 107704 380032 107710
rect 379980 107646 380032 107652
rect 379612 106956 379664 106962
rect 379612 106898 379664 106904
rect 380452 105602 380480 110092
rect 380544 110078 380834 110106
rect 380440 105596 380492 105602
rect 380440 105538 380492 105544
rect 378876 104168 378928 104174
rect 378876 104110 378928 104116
rect 380544 99374 380572 110078
rect 381188 108662 381216 110092
rect 381280 110078 381662 110106
rect 381740 110078 382030 110106
rect 382384 110078 382490 110106
rect 382568 110078 382858 110106
rect 382936 110078 383226 110106
rect 381176 108656 381228 108662
rect 381176 108598 381228 108604
rect 381280 104258 381308 110078
rect 381740 109034 381768 110078
rect 379532 99346 380572 99374
rect 380912 104230 381308 104258
rect 381464 109006 381768 109034
rect 378324 73840 378376 73846
rect 378324 73782 378376 73788
rect 379532 71058 379560 99346
rect 379520 71052 379572 71058
rect 379520 70994 379572 71000
rect 379520 53100 379572 53106
rect 379520 53042 379572 53048
rect 378324 21480 378376 21486
rect 378324 21422 378376 21428
rect 378336 16574 378364 21422
rect 378336 16546 378456 16574
rect 378232 9104 378284 9110
rect 378232 9046 378284 9052
rect 378140 4820 378192 4826
rect 378140 4762 378192 4768
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 53042
rect 380912 9042 380940 104230
rect 381464 99374 381492 109006
rect 381544 107704 381596 107710
rect 381544 107646 381596 107652
rect 381096 99346 381492 99374
rect 380992 94512 381044 94518
rect 380992 94454 381044 94460
rect 381004 16574 381032 94454
rect 381096 69698 381124 99346
rect 381556 94518 381584 107646
rect 382384 104650 382412 110078
rect 382568 109034 382596 110078
rect 382476 109006 382596 109034
rect 382372 104644 382424 104650
rect 382372 104586 382424 104592
rect 382372 104440 382424 104446
rect 382372 104382 382424 104388
rect 382280 101380 382332 101386
rect 382280 101322 382332 101328
rect 381544 94512 381596 94518
rect 381544 94454 381596 94460
rect 381084 69692 381136 69698
rect 381084 69634 381136 69640
rect 381004 16546 381216 16574
rect 380900 9036 380952 9042
rect 380900 8978 380952 8984
rect 381188 480 381216 16546
rect 382292 8974 382320 101322
rect 382384 24138 382412 104382
rect 382476 101386 382504 109006
rect 382464 101380 382516 101386
rect 382464 101322 382516 101328
rect 382936 99374 382964 110078
rect 383672 107778 383700 110092
rect 383660 107772 383712 107778
rect 383660 107714 383712 107720
rect 384040 107710 384068 110092
rect 384132 110078 384514 110106
rect 384592 110078 384882 110106
rect 385236 110078 385342 110106
rect 385420 110078 385710 110106
rect 385788 110078 386078 110106
rect 386538 110078 386644 110106
rect 384028 107704 384080 107710
rect 384028 107646 384080 107652
rect 384132 104258 384160 110078
rect 382476 99346 382964 99374
rect 383672 104230 384160 104258
rect 382476 98666 382504 99346
rect 382464 98660 382516 98666
rect 382464 98602 382516 98608
rect 382464 72480 382516 72486
rect 382464 72422 382516 72428
rect 382372 24132 382424 24138
rect 382372 24074 382424 24080
rect 382476 16574 382504 72422
rect 383672 68338 383700 104230
rect 384592 99374 384620 110078
rect 385132 104372 385184 104378
rect 385132 104314 385184 104320
rect 385040 104100 385092 104106
rect 385040 104042 385092 104048
rect 383764 99346 384620 99374
rect 383764 91798 383792 99346
rect 383752 91792 383804 91798
rect 383752 91734 383804 91740
rect 383660 68332 383712 68338
rect 383660 68274 383712 68280
rect 385052 26926 385080 104042
rect 385144 90370 385172 104314
rect 385132 90364 385184 90370
rect 385132 90306 385184 90312
rect 385236 55894 385264 110078
rect 385420 104106 385448 110078
rect 385684 107704 385736 107710
rect 385684 107646 385736 107652
rect 385408 104100 385460 104106
rect 385408 104042 385460 104048
rect 385696 57254 385724 107646
rect 385788 104378 385816 110078
rect 385868 107772 385920 107778
rect 385868 107714 385920 107720
rect 385776 104372 385828 104378
rect 385776 104314 385828 104320
rect 385880 99374 385908 107714
rect 386616 104650 386644 110078
rect 386708 110078 386906 110106
rect 386604 104644 386656 104650
rect 386604 104586 386656 104592
rect 386604 104440 386656 104446
rect 386604 104382 386656 104388
rect 386512 104100 386564 104106
rect 386512 104042 386564 104048
rect 386420 99748 386472 99754
rect 386420 99690 386472 99696
rect 385788 99346 385908 99374
rect 385788 93158 385816 99346
rect 385776 93152 385828 93158
rect 385776 93094 385828 93100
rect 385684 57248 385736 57254
rect 385684 57190 385736 57196
rect 385132 55888 385184 55894
rect 385132 55830 385184 55836
rect 385224 55888 385276 55894
rect 385224 55830 385276 55836
rect 385040 26920 385092 26926
rect 385040 26862 385092 26868
rect 383660 24200 383712 24206
rect 383660 24142 383712 24148
rect 383672 16574 383700 24142
rect 385144 16574 385172 55830
rect 386432 33794 386460 99690
rect 386524 53106 386552 104042
rect 386616 54534 386644 104382
rect 386708 99754 386736 110078
rect 387352 107710 387380 110092
rect 387444 110078 387734 110106
rect 387904 110078 388102 110106
rect 388180 110078 388562 110106
rect 388640 110078 388930 110106
rect 389192 110078 389390 110106
rect 389468 110078 389758 110106
rect 389836 110078 390126 110106
rect 387340 107704 387392 107710
rect 387340 107646 387392 107652
rect 387444 104106 387472 110078
rect 387432 104100 387484 104106
rect 387432 104042 387484 104048
rect 386696 99748 386748 99754
rect 386696 99690 386748 99696
rect 387800 89004 387852 89010
rect 387800 88946 387852 88952
rect 386696 54596 386748 54602
rect 386696 54538 386748 54544
rect 386604 54528 386656 54534
rect 386604 54470 386656 54476
rect 386512 53100 386564 53106
rect 386512 53042 386564 53048
rect 386420 33788 386472 33794
rect 386420 33730 386472 33736
rect 382476 16546 383608 16574
rect 383672 16546 384344 16574
rect 385144 16546 386000 16574
rect 382372 9444 382424 9450
rect 382372 9386 382424 9392
rect 382280 8968 382332 8974
rect 382280 8910 382332 8916
rect 382384 480 382412 9386
rect 383580 480 383608 16546
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 54538
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 88946
rect 387904 28286 387932 110078
rect 387984 104100 388036 104106
rect 387984 104042 388036 104048
rect 387996 51746 388024 104042
rect 388180 99374 388208 110078
rect 388640 104106 388668 110078
rect 388628 104100 388680 104106
rect 388628 104042 388680 104048
rect 388088 99346 388208 99374
rect 388088 89010 388116 99346
rect 388076 89004 388128 89010
rect 388076 88946 388128 88952
rect 387984 51740 388036 51746
rect 387984 51682 388036 51688
rect 389192 49026 389220 110078
rect 389272 106820 389324 106826
rect 389272 106762 389324 106768
rect 389284 50386 389312 106762
rect 389468 103514 389496 110078
rect 389836 106826 389864 110078
rect 390572 108730 390600 110092
rect 390664 110078 390954 110106
rect 391032 110078 391414 110106
rect 391492 110078 391782 110106
rect 390560 108724 390612 108730
rect 390560 108666 390612 108672
rect 389824 106820 389876 106826
rect 389824 106762 389876 106768
rect 390560 106820 390612 106826
rect 390560 106762 390612 106768
rect 389376 103486 389496 103514
rect 389376 87650 389404 103486
rect 389364 87644 389416 87650
rect 389364 87586 389416 87592
rect 389272 50380 389324 50386
rect 389272 50322 389324 50328
rect 389180 49020 389232 49026
rect 389180 48962 389232 48968
rect 389180 32428 389232 32434
rect 389180 32370 389232 32376
rect 387892 28280 387944 28286
rect 387892 28222 387944 28228
rect 389192 16574 389220 32370
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 5234 390600 106762
rect 390560 5228 390612 5234
rect 390560 5170 390612 5176
rect 390664 5114 390692 110078
rect 391032 103514 391060 110078
rect 391492 106826 391520 110078
rect 392584 108588 392636 108594
rect 392584 108530 392636 108536
rect 391480 106820 391532 106826
rect 391480 106762 391532 106768
rect 390572 5086 390692 5114
rect 390756 103486 391060 103514
rect 390572 3466 390600 5086
rect 390756 3602 390784 103486
rect 391940 93288 391992 93294
rect 391940 93230 391992 93236
rect 390836 25560 390888 25566
rect 390836 25502 390888 25508
rect 390744 3596 390796 3602
rect 390744 3538 390796 3544
rect 390848 3482 390876 25502
rect 390928 18624 390980 18630
rect 390928 18566 390980 18572
rect 390940 16574 390968 18566
rect 391952 16574 391980 93230
rect 392596 18630 392624 108530
rect 392676 107704 392728 107710
rect 392676 107646 392728 107652
rect 392688 25566 392716 107646
rect 392676 25560 392728 25566
rect 392676 25502 392728 25508
rect 393320 22772 393372 22778
rect 393320 22714 393372 22720
rect 392584 18624 392636 18630
rect 392584 18566 392636 18572
rect 393332 16574 393360 22714
rect 393976 20670 394004 119167
rect 394068 33114 394096 125423
rect 394160 60722 394188 137935
rect 394252 73166 394280 144055
rect 394344 86970 394372 150311
rect 394436 100706 394464 156567
rect 394528 113150 394556 162823
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 395344 131164 395396 131170
rect 395344 131106 395396 131112
rect 395356 115258 395384 131106
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 395344 115252 395396 115258
rect 395344 115194 395396 115200
rect 580264 115252 580316 115258
rect 580264 115194 580316 115200
rect 394516 113144 394568 113150
rect 580172 113144 580224 113150
rect 394516 113086 394568 113092
rect 394606 113112 394662 113121
rect 580172 113086 580224 113092
rect 394606 113047 394662 113056
rect 394620 111858 394648 113047
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 394608 111852 394660 111858
rect 394608 111794 394660 111800
rect 395344 111852 395396 111858
rect 395344 111794 395396 111800
rect 394424 100700 394476 100706
rect 394424 100642 394476 100648
rect 394700 100088 394752 100094
rect 394700 100030 394752 100036
rect 394332 86964 394384 86970
rect 394332 86906 394384 86912
rect 394240 73160 394292 73166
rect 394240 73102 394292 73108
rect 394148 60716 394200 60722
rect 394148 60658 394200 60664
rect 394056 33108 394108 33114
rect 394056 33050 394108 33056
rect 393964 20664 394016 20670
rect 393964 20606 394016 20612
rect 394712 16574 394740 100030
rect 395356 29646 395384 111794
rect 400864 108724 400916 108730
rect 400864 108666 400916 108672
rect 396724 108656 396776 108662
rect 396724 108598 396776 108604
rect 396080 86284 396132 86290
rect 396080 86226 396132 86232
rect 395344 29640 395396 29646
rect 395344 29582 395396 29588
rect 390940 16546 391888 16574
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390928 5228 390980 5234
rect 390928 5170 390980 5176
rect 390560 3460 390612 3466
rect 390560 3402 390612 3408
rect 390664 3454 390876 3482
rect 390664 480 390692 3454
rect 390940 3369 390968 5170
rect 390926 3360 390982 3369
rect 390926 3295 390982 3304
rect 391860 480 391888 16546
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 86226
rect 396736 22778 396764 108598
rect 398840 105732 398892 105738
rect 398840 105674 398892 105680
rect 397460 60036 397512 60042
rect 397460 59978 397512 59984
rect 396724 22772 396776 22778
rect 396724 22714 396776 22720
rect 397472 16574 397500 59978
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3074 398880 105674
rect 398932 96076 398984 96082
rect 398932 96018 398984 96024
rect 398944 3194 398972 96018
rect 400220 57316 400272 57322
rect 400220 57258 400272 57264
rect 400232 16574 400260 57258
rect 400876 47598 400904 108666
rect 429200 108520 429252 108526
rect 429200 108462 429252 108468
rect 405740 104304 405792 104310
rect 405740 104246 405792 104252
rect 402980 98796 403032 98802
rect 402980 98738 403032 98744
rect 401600 84924 401652 84930
rect 401600 84866 401652 84872
rect 400864 47592 400916 47598
rect 400864 47534 400916 47540
rect 401612 16574 401640 84866
rect 402992 16574 403020 98738
rect 404360 89072 404412 89078
rect 404360 89014 404412 89020
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 89014
rect 405752 16574 405780 104246
rect 422300 96008 422352 96014
rect 422300 95950 422352 95956
rect 418160 93220 418212 93226
rect 418160 93162 418212 93168
rect 408500 83564 408552 83570
rect 408500 83506 408552 83512
rect 407120 62892 407172 62898
rect 407120 62834 407172 62840
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3194 407160 62834
rect 408512 16574 408540 83506
rect 415400 82204 415452 82210
rect 415400 82146 415452 82152
rect 411260 29708 411312 29714
rect 411260 29650 411312 29656
rect 411272 16574 411300 29650
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 407212 10872 407264 10878
rect 407212 10814 407264 10820
rect 407120 3188 407172 3194
rect 407120 3130 407172 3136
rect 407224 480 407252 10814
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 10804 410852 10810
rect 410800 10746 410852 10752
rect 410812 480 410840 10746
rect 411916 480 411944 16546
rect 414296 10736 414348 10742
rect 414296 10678 414348 10684
rect 413100 6316 413152 6322
rect 413100 6258 413152 6264
rect 413112 480 413140 6258
rect 414308 480 414336 10678
rect 415412 3262 415440 82146
rect 415492 19984 415544 19990
rect 415492 19926 415544 19932
rect 415400 3256 415452 3262
rect 415400 3198 415452 3204
rect 415504 480 415532 19926
rect 418172 16574 418200 93162
rect 422312 16574 422340 95950
rect 426440 80776 426492 80782
rect 426440 80718 426492 80724
rect 426452 16574 426480 80718
rect 418172 16546 418568 16574
rect 422312 16546 422616 16574
rect 426452 16546 426848 16574
rect 417424 10668 417476 10674
rect 417424 10610 417476 10616
rect 416688 3256 416740 3262
rect 416688 3198 416740 3204
rect 416700 480 416728 3198
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 10610
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420920 10600 420972 10606
rect 420920 10542 420972 10548
rect 420184 6248 420236 6254
rect 420184 6190 420236 6196
rect 420196 480 420224 6190
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 10542
rect 422588 480 422616 16546
rect 423680 10532 423732 10538
rect 423680 10474 423732 10480
rect 423692 3262 423720 10474
rect 423772 6180 423824 6186
rect 423772 6122 423824 6128
rect 423680 3256 423732 3262
rect 423680 3198 423732 3204
rect 423784 480 423812 6122
rect 424968 3256 425020 3262
rect 424968 3198 425020 3204
rect 424980 480 425008 3198
rect 426164 3188 426216 3194
rect 426164 3130 426216 3136
rect 426176 480 426204 3130
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428464 10464 428516 10470
rect 428464 10406 428516 10412
rect 428476 480 428504 10406
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 108462
rect 436100 108452 436152 108458
rect 436100 108394 436152 108400
rect 430580 107092 430632 107098
rect 430580 107034 430632 107040
rect 430592 16574 430620 107034
rect 434720 91860 434772 91866
rect 434720 91802 434772 91808
rect 433340 26988 433392 26994
rect 433340 26930 433392 26936
rect 433352 16574 433380 26930
rect 434732 16574 434760 91802
rect 436112 16574 436140 108394
rect 443000 108384 443052 108390
rect 443000 108326 443052 108332
rect 441620 97368 441672 97374
rect 441620 97310 441672 97316
rect 437480 79416 437532 79422
rect 437480 79358 437532 79364
rect 430592 16546 430896 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 430868 480 430896 16546
rect 432052 10396 432104 10402
rect 432052 10338 432104 10344
rect 432064 480 432092 10338
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 79358
rect 440332 78056 440384 78062
rect 440332 77998 440384 78004
rect 439136 10328 439188 10334
rect 439136 10270 439188 10276
rect 439148 480 439176 10270
rect 440344 3398 440372 77998
rect 441632 16574 441660 97310
rect 443012 16574 443040 108326
rect 449900 108316 449952 108322
rect 449900 108258 449952 108264
rect 445760 87712 445812 87718
rect 445760 87654 445812 87660
rect 444380 76628 444432 76634
rect 444380 76570 444432 76576
rect 444392 16574 444420 76570
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 1714 440280 3334
rect 440252 1686 440372 1714
rect 440344 480 440372 1686
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 87654
rect 448520 75268 448572 75274
rect 448520 75210 448572 75216
rect 447416 4140 447468 4146
rect 447416 4082 447468 4088
rect 447428 480 447456 4082
rect 448532 3210 448560 75210
rect 448612 33856 448664 33862
rect 448612 33798 448664 33804
rect 448624 3398 448652 33798
rect 449912 16574 449940 108258
rect 480260 107024 480312 107030
rect 480260 106966 480312 106972
rect 458180 102876 458232 102882
rect 458180 102818 458232 102824
rect 456892 100020 456944 100026
rect 456892 99962 456944 99968
rect 455420 73908 455472 73914
rect 455420 73850 455472 73856
rect 452660 49088 452712 49094
rect 452660 49030 452712 49036
rect 451280 28348 451332 28354
rect 451280 28290 451332 28296
rect 451292 16574 451320 28290
rect 452672 16574 452700 49030
rect 455432 16574 455460 73850
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 454500 4072 454552 4078
rect 454500 4014 454552 4020
rect 454512 480 454540 4014
rect 455708 480 455736 16546
rect 456904 480 456932 99962
rect 458192 16574 458220 102818
rect 466460 94580 466512 94586
rect 466460 94522 466512 94528
rect 463700 90432 463752 90438
rect 463700 90374 463752 90380
rect 459560 47660 459612 47666
rect 459560 47602 459612 47608
rect 459572 16574 459600 47602
rect 463712 16574 463740 90374
rect 465172 71120 465224 71126
rect 465172 71062 465224 71068
rect 465184 16574 465212 71062
rect 466472 16574 466500 94522
rect 469220 69760 469272 69766
rect 469220 69702 469272 69708
rect 469232 16574 469260 69702
rect 470600 46232 470652 46238
rect 470600 46174 470652 46180
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 469232 16546 469904 16574
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 462780 7812 462832 7818
rect 462780 7754 462832 7760
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 462792 480 462820 7754
rect 463988 480 464016 16546
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 46174
rect 477500 44872 477552 44878
rect 477500 44814 477552 44820
rect 477512 16574 477540 44814
rect 480272 16574 480300 106966
rect 546500 106956 546552 106962
rect 546500 106898 546552 106904
rect 483020 105664 483072 105670
rect 483020 105606 483072 105612
rect 481640 68400 481692 68406
rect 481640 68342 481692 68348
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 474096 11892 474148 11898
rect 474096 11834 474148 11840
rect 473452 7744 473504 7750
rect 473452 7686 473504 7692
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 7686
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 11834
rect 476948 7676 477000 7682
rect 476948 7618 477000 7624
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 476960 480 476988 7618
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 6914 481680 68342
rect 481732 43444 481784 43450
rect 481732 43386 481784 43392
rect 481744 16574 481772 43386
rect 483032 16574 483060 105606
rect 487160 104236 487212 104242
rect 487160 104178 487212 104184
rect 484400 66904 484452 66910
rect 484400 66846 484452 66852
rect 484412 16574 484440 66846
rect 485780 42084 485832 42090
rect 485780 42026 485832 42032
rect 485792 16574 485820 42026
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 104178
rect 539600 104168 539652 104174
rect 539600 104110 539652 104116
rect 489920 102808 489972 102814
rect 489920 102750 489972 102756
rect 488540 65544 488592 65550
rect 488540 65486 488592 65492
rect 488552 16574 488580 65486
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 102750
rect 494060 101516 494112 101522
rect 494060 101458 494112 101464
rect 490012 35216 490064 35222
rect 490012 35158 490064 35164
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 35158
rect 494072 16574 494100 101458
rect 534080 101448 534132 101454
rect 534080 101390 534132 101396
rect 498200 98728 498252 98734
rect 498200 98670 498252 98676
rect 495440 84856 495492 84862
rect 495440 84798 495492 84804
rect 494072 16546 494744 16574
rect 493048 11824 493100 11830
rect 493048 11766 493100 11772
rect 492312 7608 492364 7614
rect 492312 7550 492364 7556
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 7550
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 11766
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 84798
rect 496820 36576 496872 36582
rect 496820 36518 496872 36524
rect 496832 16574 496860 36518
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 98670
rect 507860 97300 507912 97306
rect 507860 97242 507912 97248
rect 506480 83496 506532 83502
rect 506480 83438 506532 83444
rect 498292 64184 498344 64190
rect 498292 64126 498344 64132
rect 498304 16574 498332 64126
rect 502340 62824 502392 62830
rect 502340 62766 502392 62772
rect 499580 40724 499632 40730
rect 499580 40666 499632 40672
rect 499592 16574 499620 40666
rect 500960 17264 501012 17270
rect 500960 17206 501012 17212
rect 500972 16574 501000 17206
rect 502352 16574 502380 62766
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 505376 14476 505428 14482
rect 505376 14418 505428 14424
rect 503720 11756 503772 11762
rect 503720 11698 503772 11704
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 11698
rect 505388 480 505416 14418
rect 506492 480 506520 83438
rect 506572 39364 506624 39370
rect 506572 39306 506624 39312
rect 506584 16574 506612 39306
rect 507872 16574 507900 97242
rect 509240 82136 509292 82142
rect 509240 82078 509292 82084
rect 509252 16574 509280 82078
rect 520280 80708 520332 80714
rect 520280 80650 520332 80656
rect 517520 79348 517572 79354
rect 517520 79290 517572 79296
rect 513380 61396 513432 61402
rect 513380 61338 513432 61344
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 13252 511316 13258
rect 511264 13194 511316 13200
rect 511276 480 511304 13194
rect 512460 5160 512512 5166
rect 512460 5102 512512 5108
rect 512472 480 512500 5102
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 61338
rect 516140 58676 516192 58682
rect 516140 58618 516192 58624
rect 514760 37936 514812 37942
rect 514760 37878 514812 37884
rect 514772 480 514800 37878
rect 516152 16574 516180 58618
rect 517532 16574 517560 79290
rect 518900 18624 518952 18630
rect 518900 18566 518952 18572
rect 518912 16574 518940 18566
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515496 15904 515548 15910
rect 515496 15846 515548 15852
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 15846
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 80650
rect 521660 77988 521712 77994
rect 521660 77930 521712 77936
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 77930
rect 528560 76560 528612 76566
rect 528560 76502 528612 76508
rect 523040 31068 523092 31074
rect 523040 31010 523092 31016
rect 523052 3534 523080 31010
rect 523132 21412 523184 21418
rect 523132 21354 523184 21360
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 21354
rect 525432 13184 525484 13190
rect 525432 13126 525484 13132
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 13126
rect 527824 9376 527876 9382
rect 527824 9318 527876 9324
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 9318
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 76502
rect 534092 16574 534120 101390
rect 536840 95940 536892 95946
rect 536840 95882 536892 95888
rect 535460 75200 535512 75206
rect 535460 75142 535512 75148
rect 535472 16574 535500 75142
rect 536852 16574 536880 95882
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 532056 13116 532108 13122
rect 532056 13058 532108 13064
rect 531320 9308 531372 9314
rect 531320 9250 531372 9256
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 530136 480 530164 4966
rect 531332 480 531360 9250
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 13058
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 533724 480 533752 4898
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 538404 9240 538456 9246
rect 538404 9182 538456 9188
rect 538416 480 538444 9182
rect 539612 480 539640 104110
rect 542360 73840 542412 73846
rect 542360 73782 542412 73788
rect 542372 16574 542400 73782
rect 542372 16546 542768 16574
rect 541992 9172 542044 9178
rect 541992 9114 542044 9120
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 540808 480 540836 4830
rect 542004 480 542032 9114
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 545488 9104 545540 9110
rect 545488 9046 545540 9052
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 544396 480 544424 4762
rect 545500 480 545528 9046
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 106898
rect 547880 105596 547932 105602
rect 547880 105538 547932 105544
rect 547892 3534 547920 105538
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 556160 98660 556212 98666
rect 556160 98602 556212 98608
rect 547972 94512 548024 94518
rect 547972 94454 548024 94460
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547984 3346 548012 94454
rect 549260 71052 549312 71058
rect 549260 70994 549312 71000
rect 549272 16574 549300 70994
rect 553400 69692 553452 69698
rect 553400 69634 553452 69640
rect 550640 22772 550692 22778
rect 550640 22714 550692 22720
rect 550652 16574 550680 22714
rect 553412 16574 553440 69634
rect 554780 24132 554832 24138
rect 554780 24074 554832 24080
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 548708 3528 548760 3534
rect 548708 3470 548760 3476
rect 547892 3318 548012 3346
rect 547892 480 547920 3318
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3470
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 9036 552716 9042
rect 552664 8978 552716 8984
rect 552676 480 552704 8978
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 24074
rect 556172 16574 556200 98602
rect 557540 93152 557592 93158
rect 557540 93094 557592 93100
rect 557552 16574 557580 93094
rect 561680 91792 561732 91798
rect 561680 91734 561732 91740
rect 560300 68332 560352 68338
rect 560300 68274 560352 68280
rect 558920 57248 558972 57254
rect 558920 57190 558972 57196
rect 558932 16574 558960 57190
rect 560312 16574 560340 68274
rect 561692 16574 561720 91734
rect 564440 90364 564492 90370
rect 564440 90306 564492 90312
rect 563060 55888 563112 55894
rect 563060 55830 563112 55836
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 556172 480 556200 8910
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 55830
rect 564452 3534 564480 90306
rect 571984 89004 572036 89010
rect 571984 88946 572036 88952
rect 565820 54528 565872 54534
rect 565820 54470 565872 54476
rect 564532 26920 564584 26926
rect 564532 26862 564584 26868
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 26862
rect 565832 16574 565860 54470
rect 569960 53100 570012 53106
rect 569960 53042 570012 53048
rect 567200 33788 567252 33794
rect 567200 33730 567252 33736
rect 567212 16574 567240 33730
rect 568580 25560 568632 25566
rect 568580 25502 568632 25508
rect 568592 16574 568620 25502
rect 569972 16574 570000 53042
rect 570604 28280 570656 28286
rect 570604 28222 570656 28228
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 570616 3534 570644 28222
rect 571996 3534 572024 88946
rect 575480 87644 575532 87650
rect 575480 87586 575532 87592
rect 572076 51740 572128 51746
rect 572076 51682 572128 51688
rect 570604 3528 570656 3534
rect 570604 3470 570656 3476
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 571536 480 571564 3470
rect 572088 3398 572116 51682
rect 574744 50380 574796 50386
rect 574744 50322 574796 50328
rect 574100 49020 574152 49026
rect 574100 48962 574152 48968
rect 574112 16574 574140 48962
rect 574112 16546 574692 16574
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 574664 3482 574692 16546
rect 574756 3874 574784 50322
rect 575492 16574 575520 87586
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 578240 47592 578292 47598
rect 578240 47534 578292 47540
rect 578252 16574 578280 47534
rect 580276 46345 580304 115194
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580264 29640 580316 29646
rect 580264 29582 580316 29588
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 572076 3392 572128 3398
rect 572076 3334 572128 3340
rect 572732 480 572760 3470
rect 574664 3454 575152 3482
rect 573916 3392 573968 3398
rect 573916 3334 573968 3340
rect 573928 480 573956 3334
rect 575124 480 575152 3454
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 580276 6633 580304 29582
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3330 632068 3332 632088
rect 3332 632068 3384 632088
rect 3384 632068 3386 632088
rect 3330 632032 3386 632068
rect 3330 619112 3386 619168
rect 2778 606056 2834 606112
rect 3330 579944 3386 580000
rect 2962 527856 3018 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3330 501744 3386 501800
rect 3330 475632 3386 475688
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3514 658144 3570 658200
rect 3606 566888 3662 566944
rect 3422 371320 3478 371376
rect 3514 358400 3570 358456
rect 3698 553832 3754 553888
rect 3790 462576 3846 462632
rect 3606 319232 3662 319288
rect 3422 254088 3478 254144
rect 3698 306176 3754 306232
rect 3514 241032 3570 241088
rect 3422 214920 3478 214976
rect 3882 449520 3938 449576
rect 3974 423544 4030 423600
rect 3790 293120 3846 293176
rect 4066 345344 4122 345400
rect 3882 267144 3938 267200
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 189078 386552 189134 386608
rect 189078 379888 189134 379944
rect 189078 373224 189134 373280
rect 393870 368092 393872 368112
rect 393872 368092 393924 368112
rect 393924 368092 393926 368112
rect 393870 368056 393926 368092
rect 189078 366560 189134 366616
rect 394514 386824 394570 386880
rect 394606 380568 394662 380624
rect 394146 374312 394202 374368
rect 393962 361936 394018 361992
rect 189078 359896 189134 359952
rect 189078 353252 189134 353288
rect 189078 353232 189080 353252
rect 189080 353232 189132 353252
rect 189132 353232 189134 353252
rect 189078 346568 189134 346624
rect 189078 339904 189134 339960
rect 189078 333240 189134 333296
rect 393962 330792 394018 330848
rect 189078 326576 189134 326632
rect 189078 319912 189134 319968
rect 189078 313248 189134 313304
rect 189078 306584 189134 306640
rect 189078 299920 189134 299976
rect 189078 293256 189134 293312
rect 189078 286592 189134 286648
rect 393686 281016 393742 281072
rect 189078 279928 189134 279984
rect 189078 273264 189134 273320
rect 189078 266600 189134 266656
rect 189078 259936 189134 259992
rect 189078 253272 189134 253328
rect 394606 355680 394662 355736
rect 394606 349424 394662 349480
rect 394238 343168 394294 343224
rect 394606 337048 394662 337104
rect 394606 324536 394662 324592
rect 394606 318280 394662 318336
rect 394606 312160 394662 312216
rect 394238 305904 394294 305960
rect 394606 299648 394662 299704
rect 394606 293392 394662 293448
rect 394606 287272 394662 287328
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 579986 577632 580042 577688
rect 579618 537784 579674 537840
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580354 617480 580410 617536
rect 580262 378392 580318 378448
rect 580170 365064 580226 365120
rect 580170 312024 580226 312080
rect 580446 590960 580502 591016
rect 580354 351872 580410 351928
rect 394606 274760 394662 274816
rect 580262 272176 580318 272232
rect 394054 268504 394110 268560
rect 394606 262384 394662 262440
rect 580170 258848 580226 258904
rect 393962 249872 394018 249928
rect 189078 246608 189134 246664
rect 189078 239944 189134 240000
rect 189078 233280 189134 233336
rect 189078 226616 189134 226672
rect 189078 219952 189134 220008
rect 394606 256128 394662 256184
rect 394606 243616 394662 243672
rect 580538 564304 580594 564360
rect 580630 524456 580686 524512
rect 580722 511264 580778 511320
rect 580446 325216 580502 325272
rect 580814 484608 580870 484664
rect 580906 431568 580962 431624
rect 580538 298696 580594 298752
rect 580354 245520 580410 245576
rect 394606 237496 394662 237552
rect 579802 232328 579858 232384
rect 394054 231240 394110 231296
rect 394606 224984 394662 225040
rect 580170 219000 580226 219056
rect 393962 218728 394018 218784
rect 189078 213288 189134 213344
rect 393962 212608 394018 212664
rect 189078 206624 189134 206680
rect 394606 206352 394662 206408
rect 580170 205672 580226 205728
rect 3146 201864 3202 201920
rect 394054 200096 394110 200152
rect 189078 199960 189134 200016
rect 393962 193840 394018 193896
rect 189078 193296 189134 193352
rect 3422 188808 3478 188864
rect 189814 186632 189870 186688
rect 189078 179968 189134 180024
rect 3238 162832 3294 162888
rect 189722 173304 189778 173360
rect 189078 159976 189134 160032
rect 3422 149776 3478 149832
rect 3422 136720 3478 136776
rect 3330 110608 3386 110664
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 2870 32408 2926 32464
rect 189078 139984 189134 140040
rect 580170 192480 580226 192536
rect 394238 187720 394294 187776
rect 394146 181464 394202 181520
rect 394054 175208 394110 175264
rect 393962 168952 394018 169008
rect 190182 166640 190238 166696
rect 190090 153312 190146 153368
rect 189998 146648 190054 146704
rect 189906 133320 189962 133376
rect 189814 126656 189870 126712
rect 189078 119992 189134 120048
rect 189722 113328 189778 113384
rect 3606 97552 3662 97608
rect 3514 58520 3570 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 393778 131688 393834 131744
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 394514 162832 394570 162888
rect 394422 156576 394478 156632
rect 394330 150320 394386 150376
rect 394238 144064 394294 144120
rect 394146 137944 394202 138000
rect 394054 125432 394110 125488
rect 393962 119176 394018 119232
rect 193586 3576 193642 3632
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 394606 113056 394662 113112
rect 580170 112784 580226 112840
rect 390926 3304 390982 3360
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580262 6568 580318 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580349 617538 580415 617541
rect 583520 617538 584960 617628
rect 580349 617536 584960 617538
rect 580349 617480 580354 617536
rect 580410 617480 584960 617536
rect 580349 617478 584960 617480
rect 580349 617475 580415 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 579981 577690 580047 577693
rect 583520 577690 584960 577780
rect 579981 577688 584960 577690
rect 579981 577632 579986 577688
rect 580042 577632 584960 577688
rect 579981 577630 584960 577632
rect 579981 577627 580047 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 580533 564362 580599 564365
rect 583520 564362 584960 564452
rect 580533 564360 584960 564362
rect 580533 564304 580538 564360
rect 580594 564304 584960 564360
rect 580533 564302 584960 564304
rect 580533 564299 580599 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579613 537842 579679 537845
rect 583520 537842 584960 537932
rect 579613 537840 584960 537842
rect 579613 537784 579618 537840
rect 579674 537784 584960 537840
rect 579613 537782 584960 537784
rect 579613 537779 579679 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580625 524514 580691 524517
rect 583520 524514 584960 524604
rect 580625 524512 584960 524514
rect 580625 524456 580630 524512
rect 580686 524456 584960 524512
rect 580625 524454 584960 524456
rect 580625 524451 580691 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580717 511322 580783 511325
rect 583520 511322 584960 511412
rect 580717 511320 584960 511322
rect 580717 511264 580722 511320
rect 580778 511264 584960 511320
rect 580717 511262 584960 511264
rect 580717 511259 580783 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580809 484666 580875 484669
rect 583520 484666 584960 484756
rect 580809 484664 584960 484666
rect 580809 484608 580814 484664
rect 580870 484608 584960 484664
rect 580809 484606 584960 484608
rect 580809 484603 580875 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3785 462634 3851 462637
rect -960 462632 3851 462634
rect -960 462576 3790 462632
rect 3846 462576 3851 462632
rect -960 462574 3851 462576
rect -960 462484 480 462574
rect 3785 462571 3851 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3877 449578 3943 449581
rect -960 449576 3943 449578
rect -960 449520 3882 449576
rect 3938 449520 3943 449576
rect -960 449518 3943 449520
rect -960 449428 480 449518
rect 3877 449515 3943 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3969 423602 4035 423605
rect -960 423600 4035 423602
rect -960 423544 3974 423600
rect 4030 423544 4035 423600
rect -960 423542 4035 423544
rect -960 423452 480 423542
rect 3969 423539 4035 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect 394509 386882 394575 386885
rect 391828 386880 394575 386882
rect 391828 386824 394514 386880
rect 394570 386824 394575 386880
rect 391828 386822 394575 386824
rect 394509 386819 394575 386822
rect 189073 386610 189139 386613
rect 189073 386608 192188 386610
rect 189073 386552 189078 386608
rect 189134 386552 192188 386608
rect 189073 386550 192188 386552
rect 189073 386547 189139 386550
rect -960 384284 480 384524
rect 394601 380626 394667 380629
rect 391828 380624 394667 380626
rect 391828 380568 394606 380624
rect 394662 380568 394667 380624
rect 391828 380566 394667 380568
rect 394601 380563 394667 380566
rect 189073 379946 189139 379949
rect 189073 379944 192188 379946
rect 189073 379888 189078 379944
rect 189134 379888 192188 379944
rect 189073 379886 192188 379888
rect 189073 379883 189139 379886
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 394141 374370 394207 374373
rect 391828 374368 394207 374370
rect 391828 374312 394146 374368
rect 394202 374312 394207 374368
rect 391828 374310 394207 374312
rect 394141 374307 394207 374310
rect 189073 373282 189139 373285
rect 189073 373280 192188 373282
rect 189073 373224 189078 373280
rect 189134 373224 192188 373280
rect 189073 373222 192188 373224
rect 189073 373219 189139 373222
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 393865 368114 393931 368117
rect 391828 368112 393931 368114
rect 391828 368056 393870 368112
rect 393926 368056 393931 368112
rect 391828 368054 393931 368056
rect 393865 368051 393931 368054
rect 189073 366618 189139 366621
rect 189073 366616 192188 366618
rect 189073 366560 189078 366616
rect 189134 366560 192188 366616
rect 189073 366558 192188 366560
rect 189073 366555 189139 366558
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 393957 361994 394023 361997
rect 391828 361992 394023 361994
rect 391828 361936 393962 361992
rect 394018 361936 394023 361992
rect 391828 361934 394023 361936
rect 393957 361931 394023 361934
rect 189073 359954 189139 359957
rect 189073 359952 192188 359954
rect 189073 359896 189078 359952
rect 189134 359896 192188 359952
rect 189073 359894 192188 359896
rect 189073 359891 189139 359894
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 394601 355738 394667 355741
rect 391828 355736 394667 355738
rect 391828 355680 394606 355736
rect 394662 355680 394667 355736
rect 391828 355678 394667 355680
rect 394601 355675 394667 355678
rect 189073 353290 189139 353293
rect 189073 353288 192188 353290
rect 189073 353232 189078 353288
rect 189134 353232 192188 353288
rect 189073 353230 192188 353232
rect 189073 353227 189139 353230
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 394601 349482 394667 349485
rect 391828 349480 394667 349482
rect 391828 349424 394606 349480
rect 394662 349424 394667 349480
rect 391828 349422 394667 349424
rect 394601 349419 394667 349422
rect 189073 346626 189139 346629
rect 189073 346624 192188 346626
rect 189073 346568 189078 346624
rect 189134 346568 192188 346624
rect 189073 346566 192188 346568
rect 189073 346563 189139 346566
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 394233 343226 394299 343229
rect 391828 343224 394299 343226
rect 391828 343168 394238 343224
rect 394294 343168 394299 343224
rect 391828 343166 394299 343168
rect 394233 343163 394299 343166
rect 189073 339962 189139 339965
rect 189073 339960 192188 339962
rect 189073 339904 189078 339960
rect 189134 339904 192188 339960
rect 189073 339902 192188 339904
rect 189073 339899 189139 339902
rect 583520 338452 584960 338692
rect 394601 337106 394667 337109
rect 391828 337104 394667 337106
rect 391828 337048 394606 337104
rect 394662 337048 394667 337104
rect 391828 337046 394667 337048
rect 394601 337043 394667 337046
rect 189073 333298 189139 333301
rect 189073 333296 192188 333298
rect 189073 333240 189078 333296
rect 189134 333240 192188 333296
rect 189073 333238 192188 333240
rect 189073 333235 189139 333238
rect -960 332196 480 332436
rect 393957 330850 394023 330853
rect 391828 330848 394023 330850
rect 391828 330792 393962 330848
rect 394018 330792 394023 330848
rect 391828 330790 394023 330792
rect 393957 330787 394023 330790
rect 189073 326634 189139 326637
rect 189073 326632 192188 326634
rect 189073 326576 189078 326632
rect 189134 326576 192188 326632
rect 189073 326574 192188 326576
rect 189073 326571 189139 326574
rect 580441 325274 580507 325277
rect 583520 325274 584960 325364
rect 580441 325272 584960 325274
rect 580441 325216 580446 325272
rect 580502 325216 584960 325272
rect 580441 325214 584960 325216
rect 580441 325211 580507 325214
rect 583520 325124 584960 325214
rect 394601 324594 394667 324597
rect 391828 324592 394667 324594
rect 391828 324536 394606 324592
rect 394662 324536 394667 324592
rect 391828 324534 394667 324536
rect 394601 324531 394667 324534
rect 189073 319970 189139 319973
rect 189073 319968 192188 319970
rect 189073 319912 189078 319968
rect 189134 319912 192188 319968
rect 189073 319910 192188 319912
rect 189073 319907 189139 319910
rect -960 319290 480 319380
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 394601 318338 394667 318341
rect 391828 318336 394667 318338
rect 391828 318280 394606 318336
rect 394662 318280 394667 318336
rect 391828 318278 394667 318280
rect 394601 318275 394667 318278
rect 189073 313306 189139 313309
rect 189073 313304 192188 313306
rect 189073 313248 189078 313304
rect 189134 313248 192188 313304
rect 189073 313246 192188 313248
rect 189073 313243 189139 313246
rect 394601 312218 394667 312221
rect 391828 312216 394667 312218
rect 391828 312160 394606 312216
rect 394662 312160 394667 312216
rect 391828 312158 394667 312160
rect 394601 312155 394667 312158
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 189073 306642 189139 306645
rect 189073 306640 192188 306642
rect 189073 306584 189078 306640
rect 189134 306584 192188 306640
rect 189073 306582 192188 306584
rect 189073 306579 189139 306582
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 394233 305962 394299 305965
rect 391828 305960 394299 305962
rect 391828 305904 394238 305960
rect 394294 305904 394299 305960
rect 391828 305902 394299 305904
rect 394233 305899 394299 305902
rect 189073 299978 189139 299981
rect 189073 299976 192188 299978
rect 189073 299920 189078 299976
rect 189134 299920 192188 299976
rect 189073 299918 192188 299920
rect 189073 299915 189139 299918
rect 394601 299706 394667 299709
rect 391828 299704 394667 299706
rect 391828 299648 394606 299704
rect 394662 299648 394667 299704
rect 391828 299646 394667 299648
rect 394601 299643 394667 299646
rect 580533 298754 580599 298757
rect 583520 298754 584960 298844
rect 580533 298752 584960 298754
rect 580533 298696 580538 298752
rect 580594 298696 584960 298752
rect 580533 298694 584960 298696
rect 580533 298691 580599 298694
rect 583520 298604 584960 298694
rect 394601 293450 394667 293453
rect 391828 293448 394667 293450
rect 391828 293392 394606 293448
rect 394662 293392 394667 293448
rect 391828 293390 394667 293392
rect 394601 293387 394667 293390
rect 189073 293314 189139 293317
rect 189073 293312 192188 293314
rect -960 293178 480 293268
rect 189073 293256 189078 293312
rect 189134 293256 192188 293312
rect 189073 293254 192188 293256
rect 189073 293251 189139 293254
rect 3785 293178 3851 293181
rect -960 293176 3851 293178
rect -960 293120 3790 293176
rect 3846 293120 3851 293176
rect -960 293118 3851 293120
rect -960 293028 480 293118
rect 3785 293115 3851 293118
rect 394601 287330 394667 287333
rect 391828 287328 394667 287330
rect 391828 287272 394606 287328
rect 394662 287272 394667 287328
rect 391828 287270 394667 287272
rect 394601 287267 394667 287270
rect 189073 286650 189139 286653
rect 189073 286648 192188 286650
rect 189073 286592 189078 286648
rect 189134 286592 192188 286648
rect 189073 286590 192188 286592
rect 189073 286587 189139 286590
rect 583520 285276 584960 285516
rect 393681 281074 393747 281077
rect 391828 281072 393747 281074
rect 391828 281016 393686 281072
rect 393742 281016 393747 281072
rect 391828 281014 393747 281016
rect 393681 281011 393747 281014
rect -960 279972 480 280212
rect 189073 279986 189139 279989
rect 189073 279984 192188 279986
rect 189073 279928 189078 279984
rect 189134 279928 192188 279984
rect 189073 279926 192188 279928
rect 189073 279923 189139 279926
rect 394601 274818 394667 274821
rect 391828 274816 394667 274818
rect 391828 274760 394606 274816
rect 394662 274760 394667 274816
rect 391828 274758 394667 274760
rect 394601 274755 394667 274758
rect 189073 273322 189139 273325
rect 189073 273320 192188 273322
rect 189073 273264 189078 273320
rect 189134 273264 192188 273320
rect 189073 273262 192188 273264
rect 189073 273259 189139 273262
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 583520 272084 584960 272174
rect 394049 268562 394115 268565
rect 391828 268560 394115 268562
rect 391828 268504 394054 268560
rect 394110 268504 394115 268560
rect 391828 268502 394115 268504
rect 394049 268499 394115 268502
rect -960 267202 480 267292
rect 3877 267202 3943 267205
rect -960 267200 3943 267202
rect -960 267144 3882 267200
rect 3938 267144 3943 267200
rect -960 267142 3943 267144
rect -960 267052 480 267142
rect 3877 267139 3943 267142
rect 189073 266658 189139 266661
rect 189073 266656 192188 266658
rect 189073 266600 189078 266656
rect 189134 266600 192188 266656
rect 189073 266598 192188 266600
rect 189073 266595 189139 266598
rect 394601 262442 394667 262445
rect 391828 262440 394667 262442
rect 391828 262384 394606 262440
rect 394662 262384 394667 262440
rect 391828 262382 394667 262384
rect 394601 262379 394667 262382
rect 189073 259994 189139 259997
rect 189073 259992 192188 259994
rect 189073 259936 189078 259992
rect 189134 259936 192188 259992
rect 189073 259934 192188 259936
rect 189073 259931 189139 259934
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 394601 256186 394667 256189
rect 391828 256184 394667 256186
rect 391828 256128 394606 256184
rect 394662 256128 394667 256184
rect 391828 256126 394667 256128
rect 394601 256123 394667 256126
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 189073 253330 189139 253333
rect 189073 253328 192188 253330
rect 189073 253272 189078 253328
rect 189134 253272 192188 253328
rect 189073 253270 192188 253272
rect 189073 253267 189139 253270
rect 393957 249930 394023 249933
rect 391828 249928 394023 249930
rect 391828 249872 393962 249928
rect 394018 249872 394023 249928
rect 391828 249870 394023 249872
rect 393957 249867 394023 249870
rect 189073 246666 189139 246669
rect 189073 246664 192188 246666
rect 189073 246608 189078 246664
rect 189134 246608 192188 246664
rect 189073 246606 192188 246608
rect 189073 246603 189139 246606
rect 580349 245578 580415 245581
rect 583520 245578 584960 245668
rect 580349 245576 584960 245578
rect 580349 245520 580354 245576
rect 580410 245520 584960 245576
rect 580349 245518 584960 245520
rect 580349 245515 580415 245518
rect 583520 245428 584960 245518
rect 394601 243674 394667 243677
rect 391828 243672 394667 243674
rect 391828 243616 394606 243672
rect 394662 243616 394667 243672
rect 391828 243614 394667 243616
rect 394601 243611 394667 243614
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 189073 240002 189139 240005
rect 189073 240000 192188 240002
rect 189073 239944 189078 240000
rect 189134 239944 192188 240000
rect 189073 239942 192188 239944
rect 189073 239939 189139 239942
rect 394601 237554 394667 237557
rect 391828 237552 394667 237554
rect 391828 237496 394606 237552
rect 394662 237496 394667 237552
rect 391828 237494 394667 237496
rect 394601 237491 394667 237494
rect 189073 233338 189139 233341
rect 189073 233336 192188 233338
rect 189073 233280 189078 233336
rect 189134 233280 192188 233336
rect 189073 233278 192188 233280
rect 189073 233275 189139 233278
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect 394049 231298 394115 231301
rect 391828 231296 394115 231298
rect 391828 231240 394054 231296
rect 394110 231240 394115 231296
rect 391828 231238 394115 231240
rect 394049 231235 394115 231238
rect -960 227884 480 228124
rect 189073 226674 189139 226677
rect 189073 226672 192188 226674
rect 189073 226616 189078 226672
rect 189134 226616 192188 226672
rect 189073 226614 192188 226616
rect 189073 226611 189139 226614
rect 394601 225042 394667 225045
rect 391828 225040 394667 225042
rect 391828 224984 394606 225040
rect 394662 224984 394667 225040
rect 391828 224982 394667 224984
rect 394601 224979 394667 224982
rect 189073 220010 189139 220013
rect 189073 220008 192188 220010
rect 189073 219952 189078 220008
rect 189134 219952 192188 220008
rect 189073 219950 192188 219952
rect 189073 219947 189139 219950
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 393957 218786 394023 218789
rect 391828 218784 394023 218786
rect 391828 218728 393962 218784
rect 394018 218728 394023 218784
rect 391828 218726 394023 218728
rect 393957 218723 394023 218726
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 189073 213346 189139 213349
rect 189073 213344 192188 213346
rect 189073 213288 189078 213344
rect 189134 213288 192188 213344
rect 189073 213286 192188 213288
rect 189073 213283 189139 213286
rect 393957 212666 394023 212669
rect 391828 212664 394023 212666
rect 391828 212608 393962 212664
rect 394018 212608 394023 212664
rect 391828 212606 394023 212608
rect 393957 212603 394023 212606
rect 189073 206682 189139 206685
rect 189073 206680 192188 206682
rect 189073 206624 189078 206680
rect 189134 206624 192188 206680
rect 189073 206622 192188 206624
rect 189073 206619 189139 206622
rect 394601 206410 394667 206413
rect 391828 206408 394667 206410
rect 391828 206352 394606 206408
rect 394662 206352 394667 206408
rect 391828 206350 394667 206352
rect 394601 206347 394667 206350
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3141 201922 3207 201925
rect -960 201920 3207 201922
rect -960 201864 3146 201920
rect 3202 201864 3207 201920
rect -960 201862 3207 201864
rect -960 201772 480 201862
rect 3141 201859 3207 201862
rect 394049 200154 394115 200157
rect 391828 200152 394115 200154
rect 391828 200096 394054 200152
rect 394110 200096 394115 200152
rect 391828 200094 394115 200096
rect 394049 200091 394115 200094
rect 189073 200018 189139 200021
rect 189073 200016 192188 200018
rect 189073 199960 189078 200016
rect 189134 199960 192188 200016
rect 189073 199958 192188 199960
rect 189073 199955 189139 199958
rect 393957 193898 394023 193901
rect 391828 193896 394023 193898
rect 391828 193840 393962 193896
rect 394018 193840 394023 193896
rect 391828 193838 394023 193840
rect 393957 193835 394023 193838
rect 189073 193354 189139 193357
rect 189073 193352 192188 193354
rect 189073 193296 189078 193352
rect 189134 193296 192188 193352
rect 189073 193294 192188 193296
rect 189073 193291 189139 193294
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 394233 187778 394299 187781
rect 391828 187776 394299 187778
rect 391828 187720 394238 187776
rect 394294 187720 394299 187776
rect 391828 187718 394299 187720
rect 394233 187715 394299 187718
rect 189809 186690 189875 186693
rect 189809 186688 192188 186690
rect 189809 186632 189814 186688
rect 189870 186632 192188 186688
rect 189809 186630 192188 186632
rect 189809 186627 189875 186630
rect 394141 181522 394207 181525
rect 391828 181520 394207 181522
rect 391828 181464 394146 181520
rect 394202 181464 394207 181520
rect 391828 181462 394207 181464
rect 394141 181459 394207 181462
rect 189073 180026 189139 180029
rect 189073 180024 192188 180026
rect 189073 179968 189078 180024
rect 189134 179968 192188 180024
rect 189073 179966 192188 179968
rect 189073 179963 189139 179966
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 394049 175266 394115 175269
rect 391828 175264 394115 175266
rect 391828 175208 394054 175264
rect 394110 175208 394115 175264
rect 391828 175206 394115 175208
rect 394049 175203 394115 175206
rect 189717 173362 189783 173365
rect 189717 173360 192188 173362
rect 189717 173304 189722 173360
rect 189778 173304 192188 173360
rect 189717 173302 192188 173304
rect 189717 173299 189783 173302
rect 393957 169010 394023 169013
rect 391828 169008 394023 169010
rect 391828 168952 393962 169008
rect 394018 168952 394023 169008
rect 391828 168950 394023 168952
rect 393957 168947 394023 168950
rect 190177 166698 190243 166701
rect 190177 166696 192188 166698
rect 190177 166640 190182 166696
rect 190238 166640 192188 166696
rect 190177 166638 192188 166640
rect 190177 166635 190243 166638
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect 394509 162890 394575 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 391828 162888 394575 162890
rect 391828 162832 394514 162888
rect 394570 162832 394575 162888
rect 391828 162830 394575 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 394509 162827 394575 162830
rect 189073 160034 189139 160037
rect 189073 160032 192188 160034
rect 189073 159976 189078 160032
rect 189134 159976 192188 160032
rect 189073 159974 192188 159976
rect 189073 159971 189139 159974
rect 394417 156634 394483 156637
rect 391828 156632 394483 156634
rect 391828 156576 394422 156632
rect 394478 156576 394483 156632
rect 391828 156574 394483 156576
rect 394417 156571 394483 156574
rect 190085 153370 190151 153373
rect 190085 153368 192188 153370
rect 190085 153312 190090 153368
rect 190146 153312 192188 153368
rect 190085 153310 192188 153312
rect 190085 153307 190151 153310
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 394325 150378 394391 150381
rect 391828 150376 394391 150378
rect 391828 150320 394330 150376
rect 394386 150320 394391 150376
rect 391828 150318 394391 150320
rect 394325 150315 394391 150318
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 189993 146706 190059 146709
rect 189993 146704 192188 146706
rect 189993 146648 189998 146704
rect 190054 146648 192188 146704
rect 189993 146646 192188 146648
rect 189993 146643 190059 146646
rect 394233 144122 394299 144125
rect 391828 144120 394299 144122
rect 391828 144064 394238 144120
rect 394294 144064 394299 144120
rect 391828 144062 394299 144064
rect 394233 144059 394299 144062
rect 189073 140042 189139 140045
rect 189073 140040 192188 140042
rect 189073 139984 189078 140040
rect 189134 139984 192188 140040
rect 189073 139982 192188 139984
rect 189073 139979 189139 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 394141 138002 394207 138005
rect 391828 138000 394207 138002
rect 391828 137944 394146 138000
rect 394202 137944 394207 138000
rect 391828 137942 394207 137944
rect 394141 137939 394207 137942
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 189901 133378 189967 133381
rect 189901 133376 192188 133378
rect 189901 133320 189906 133376
rect 189962 133320 192188 133376
rect 189901 133318 192188 133320
rect 189901 133315 189967 133318
rect 393773 131746 393839 131749
rect 391828 131744 393839 131746
rect 391828 131688 393778 131744
rect 393834 131688 393839 131744
rect 391828 131686 393839 131688
rect 393773 131683 393839 131686
rect 189809 126714 189875 126717
rect 189809 126712 192188 126714
rect 189809 126656 189814 126712
rect 189870 126656 192188 126712
rect 189809 126654 192188 126656
rect 189809 126651 189875 126654
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 394049 125490 394115 125493
rect 391828 125488 394115 125490
rect 391828 125432 394054 125488
rect 394110 125432 394115 125488
rect 391828 125430 394115 125432
rect 394049 125427 394115 125430
rect -960 123572 480 123812
rect 189073 120050 189139 120053
rect 189073 120048 192188 120050
rect 189073 119992 189078 120048
rect 189134 119992 192188 120048
rect 189073 119990 192188 119992
rect 189073 119987 189139 119990
rect 393957 119234 394023 119237
rect 391828 119232 394023 119234
rect 391828 119176 393962 119232
rect 394018 119176 394023 119232
rect 391828 119174 394023 119176
rect 393957 119171 394023 119174
rect 189717 113386 189783 113389
rect 189717 113384 192188 113386
rect 189717 113328 189722 113384
rect 189778 113328 192188 113384
rect 189717 113326 192188 113328
rect 189717 113323 189783 113326
rect 394601 113114 394667 113117
rect 391828 113112 394667 113114
rect 391828 113056 394606 113112
rect 394662 113056 394667 113112
rect 391828 113054 394667 113056
rect 394601 113051 394667 113054
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 193581 3634 193647 3637
rect 180750 3632 193647 3634
rect 180750 3576 193586 3632
rect 193642 3576 193647 3632
rect 180750 3574 193647 3576
rect 5257 3362 5323 3365
rect 180750 3362 180810 3574
rect 193581 3571 193647 3574
rect 5257 3360 180810 3362
rect 5257 3304 5262 3360
rect 5318 3304 180810 3360
rect 5257 3302 180810 3304
rect 390921 3362 390987 3365
rect 583385 3362 583451 3365
rect 390921 3360 583451 3362
rect 390921 3304 390926 3360
rect 390982 3304 583390 3360
rect 583446 3304 583451 3360
rect 390921 3302 583451 3304
rect 5257 3299 5323 3302
rect 390921 3299 390987 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 392000 191414 407898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 392000 195914 412398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 392000 200414 416898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 392000 204914 421398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 392000 209414 425898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 392000 213914 394398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 392000 218414 398898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 392000 222914 403398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 392000 227414 407898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 392000 231914 412398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 392000 236414 416898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 392000 240914 421398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 392000 245414 425898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 392000 249914 394398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 392000 254414 398898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 392000 258914 403398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 392000 263414 407898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 392000 267914 412398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 392000 272414 416898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 392000 276914 421398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 392000 281414 425898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 392000 285914 394398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 392000 290414 398898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 392000 294914 403398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 392000 299414 407898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 392000 303914 412398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 392000 308414 416898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 392000 312914 421398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 392000 317414 425898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 392000 321914 394398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 392000 326414 398898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 392000 330914 403398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 392000 335414 407898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 392000 339914 412398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 392000 344414 416898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 392000 348914 421398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 392000 353414 425898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 392000 357914 394398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 392000 362414 398898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 392000 366914 403398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 392000 371414 407898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 392000 375914 412398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 392000 380414 416898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 392000 384914 421398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 392000 389414 425898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 392000 393914 394398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 211568 367954 211888 367986
rect 211568 367718 211610 367954
rect 211846 367718 211888 367954
rect 211568 367634 211888 367718
rect 211568 367398 211610 367634
rect 211846 367398 211888 367634
rect 211568 367366 211888 367398
rect 242288 367954 242608 367986
rect 242288 367718 242330 367954
rect 242566 367718 242608 367954
rect 242288 367634 242608 367718
rect 242288 367398 242330 367634
rect 242566 367398 242608 367634
rect 242288 367366 242608 367398
rect 273008 367954 273328 367986
rect 273008 367718 273050 367954
rect 273286 367718 273328 367954
rect 273008 367634 273328 367718
rect 273008 367398 273050 367634
rect 273286 367398 273328 367634
rect 273008 367366 273328 367398
rect 303728 367954 304048 367986
rect 303728 367718 303770 367954
rect 304006 367718 304048 367954
rect 303728 367634 304048 367718
rect 303728 367398 303770 367634
rect 304006 367398 304048 367634
rect 303728 367366 304048 367398
rect 334448 367954 334768 367986
rect 334448 367718 334490 367954
rect 334726 367718 334768 367954
rect 334448 367634 334768 367718
rect 334448 367398 334490 367634
rect 334726 367398 334768 367634
rect 334448 367366 334768 367398
rect 365168 367954 365488 367986
rect 365168 367718 365210 367954
rect 365446 367718 365488 367954
rect 365168 367634 365488 367718
rect 365168 367398 365210 367634
rect 365446 367398 365488 367634
rect 365168 367366 365488 367398
rect 196208 363454 196528 363486
rect 196208 363218 196250 363454
rect 196486 363218 196528 363454
rect 196208 363134 196528 363218
rect 196208 362898 196250 363134
rect 196486 362898 196528 363134
rect 196208 362866 196528 362898
rect 226928 363454 227248 363486
rect 226928 363218 226970 363454
rect 227206 363218 227248 363454
rect 226928 363134 227248 363218
rect 226928 362898 226970 363134
rect 227206 362898 227248 363134
rect 226928 362866 227248 362898
rect 257648 363454 257968 363486
rect 257648 363218 257690 363454
rect 257926 363218 257968 363454
rect 257648 363134 257968 363218
rect 257648 362898 257690 363134
rect 257926 362898 257968 363134
rect 257648 362866 257968 362898
rect 288368 363454 288688 363486
rect 288368 363218 288410 363454
rect 288646 363218 288688 363454
rect 288368 363134 288688 363218
rect 288368 362898 288410 363134
rect 288646 362898 288688 363134
rect 288368 362866 288688 362898
rect 319088 363454 319408 363486
rect 319088 363218 319130 363454
rect 319366 363218 319408 363454
rect 319088 363134 319408 363218
rect 319088 362898 319130 363134
rect 319366 362898 319408 363134
rect 319088 362866 319408 362898
rect 349808 363454 350128 363486
rect 349808 363218 349850 363454
rect 350086 363218 350128 363454
rect 349808 363134 350128 363218
rect 349808 362898 349850 363134
rect 350086 362898 350128 363134
rect 349808 362866 350128 362898
rect 380528 363454 380848 363486
rect 380528 363218 380570 363454
rect 380806 363218 380848 363454
rect 380528 363134 380848 363218
rect 380528 362898 380570 363134
rect 380806 362898 380848 363134
rect 380528 362866 380848 362898
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 211568 331954 211888 331986
rect 211568 331718 211610 331954
rect 211846 331718 211888 331954
rect 211568 331634 211888 331718
rect 211568 331398 211610 331634
rect 211846 331398 211888 331634
rect 211568 331366 211888 331398
rect 242288 331954 242608 331986
rect 242288 331718 242330 331954
rect 242566 331718 242608 331954
rect 242288 331634 242608 331718
rect 242288 331398 242330 331634
rect 242566 331398 242608 331634
rect 242288 331366 242608 331398
rect 273008 331954 273328 331986
rect 273008 331718 273050 331954
rect 273286 331718 273328 331954
rect 273008 331634 273328 331718
rect 273008 331398 273050 331634
rect 273286 331398 273328 331634
rect 273008 331366 273328 331398
rect 303728 331954 304048 331986
rect 303728 331718 303770 331954
rect 304006 331718 304048 331954
rect 303728 331634 304048 331718
rect 303728 331398 303770 331634
rect 304006 331398 304048 331634
rect 303728 331366 304048 331398
rect 334448 331954 334768 331986
rect 334448 331718 334490 331954
rect 334726 331718 334768 331954
rect 334448 331634 334768 331718
rect 334448 331398 334490 331634
rect 334726 331398 334768 331634
rect 334448 331366 334768 331398
rect 365168 331954 365488 331986
rect 365168 331718 365210 331954
rect 365446 331718 365488 331954
rect 365168 331634 365488 331718
rect 365168 331398 365210 331634
rect 365446 331398 365488 331634
rect 365168 331366 365488 331398
rect 196208 327454 196528 327486
rect 196208 327218 196250 327454
rect 196486 327218 196528 327454
rect 196208 327134 196528 327218
rect 196208 326898 196250 327134
rect 196486 326898 196528 327134
rect 196208 326866 196528 326898
rect 226928 327454 227248 327486
rect 226928 327218 226970 327454
rect 227206 327218 227248 327454
rect 226928 327134 227248 327218
rect 226928 326898 226970 327134
rect 227206 326898 227248 327134
rect 226928 326866 227248 326898
rect 257648 327454 257968 327486
rect 257648 327218 257690 327454
rect 257926 327218 257968 327454
rect 257648 327134 257968 327218
rect 257648 326898 257690 327134
rect 257926 326898 257968 327134
rect 257648 326866 257968 326898
rect 288368 327454 288688 327486
rect 288368 327218 288410 327454
rect 288646 327218 288688 327454
rect 288368 327134 288688 327218
rect 288368 326898 288410 327134
rect 288646 326898 288688 327134
rect 288368 326866 288688 326898
rect 319088 327454 319408 327486
rect 319088 327218 319130 327454
rect 319366 327218 319408 327454
rect 319088 327134 319408 327218
rect 319088 326898 319130 327134
rect 319366 326898 319408 327134
rect 319088 326866 319408 326898
rect 349808 327454 350128 327486
rect 349808 327218 349850 327454
rect 350086 327218 350128 327454
rect 349808 327134 350128 327218
rect 349808 326898 349850 327134
rect 350086 326898 350128 327134
rect 349808 326866 350128 326898
rect 380528 327454 380848 327486
rect 380528 327218 380570 327454
rect 380806 327218 380848 327454
rect 380528 327134 380848 327218
rect 380528 326898 380570 327134
rect 380806 326898 380848 327134
rect 380528 326866 380848 326898
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 211568 295954 211888 295986
rect 211568 295718 211610 295954
rect 211846 295718 211888 295954
rect 211568 295634 211888 295718
rect 211568 295398 211610 295634
rect 211846 295398 211888 295634
rect 211568 295366 211888 295398
rect 242288 295954 242608 295986
rect 242288 295718 242330 295954
rect 242566 295718 242608 295954
rect 242288 295634 242608 295718
rect 242288 295398 242330 295634
rect 242566 295398 242608 295634
rect 242288 295366 242608 295398
rect 273008 295954 273328 295986
rect 273008 295718 273050 295954
rect 273286 295718 273328 295954
rect 273008 295634 273328 295718
rect 273008 295398 273050 295634
rect 273286 295398 273328 295634
rect 273008 295366 273328 295398
rect 303728 295954 304048 295986
rect 303728 295718 303770 295954
rect 304006 295718 304048 295954
rect 303728 295634 304048 295718
rect 303728 295398 303770 295634
rect 304006 295398 304048 295634
rect 303728 295366 304048 295398
rect 334448 295954 334768 295986
rect 334448 295718 334490 295954
rect 334726 295718 334768 295954
rect 334448 295634 334768 295718
rect 334448 295398 334490 295634
rect 334726 295398 334768 295634
rect 334448 295366 334768 295398
rect 365168 295954 365488 295986
rect 365168 295718 365210 295954
rect 365446 295718 365488 295954
rect 365168 295634 365488 295718
rect 365168 295398 365210 295634
rect 365446 295398 365488 295634
rect 365168 295366 365488 295398
rect 196208 291454 196528 291486
rect 196208 291218 196250 291454
rect 196486 291218 196528 291454
rect 196208 291134 196528 291218
rect 196208 290898 196250 291134
rect 196486 290898 196528 291134
rect 196208 290866 196528 290898
rect 226928 291454 227248 291486
rect 226928 291218 226970 291454
rect 227206 291218 227248 291454
rect 226928 291134 227248 291218
rect 226928 290898 226970 291134
rect 227206 290898 227248 291134
rect 226928 290866 227248 290898
rect 257648 291454 257968 291486
rect 257648 291218 257690 291454
rect 257926 291218 257968 291454
rect 257648 291134 257968 291218
rect 257648 290898 257690 291134
rect 257926 290898 257968 291134
rect 257648 290866 257968 290898
rect 288368 291454 288688 291486
rect 288368 291218 288410 291454
rect 288646 291218 288688 291454
rect 288368 291134 288688 291218
rect 288368 290898 288410 291134
rect 288646 290898 288688 291134
rect 288368 290866 288688 290898
rect 319088 291454 319408 291486
rect 319088 291218 319130 291454
rect 319366 291218 319408 291454
rect 319088 291134 319408 291218
rect 319088 290898 319130 291134
rect 319366 290898 319408 291134
rect 319088 290866 319408 290898
rect 349808 291454 350128 291486
rect 349808 291218 349850 291454
rect 350086 291218 350128 291454
rect 349808 291134 350128 291218
rect 349808 290898 349850 291134
rect 350086 290898 350128 291134
rect 349808 290866 350128 290898
rect 380528 291454 380848 291486
rect 380528 291218 380570 291454
rect 380806 291218 380848 291454
rect 380528 291134 380848 291218
rect 380528 290898 380570 291134
rect 380806 290898 380848 291134
rect 380528 290866 380848 290898
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 211568 259954 211888 259986
rect 211568 259718 211610 259954
rect 211846 259718 211888 259954
rect 211568 259634 211888 259718
rect 211568 259398 211610 259634
rect 211846 259398 211888 259634
rect 211568 259366 211888 259398
rect 242288 259954 242608 259986
rect 242288 259718 242330 259954
rect 242566 259718 242608 259954
rect 242288 259634 242608 259718
rect 242288 259398 242330 259634
rect 242566 259398 242608 259634
rect 242288 259366 242608 259398
rect 273008 259954 273328 259986
rect 273008 259718 273050 259954
rect 273286 259718 273328 259954
rect 273008 259634 273328 259718
rect 273008 259398 273050 259634
rect 273286 259398 273328 259634
rect 273008 259366 273328 259398
rect 303728 259954 304048 259986
rect 303728 259718 303770 259954
rect 304006 259718 304048 259954
rect 303728 259634 304048 259718
rect 303728 259398 303770 259634
rect 304006 259398 304048 259634
rect 303728 259366 304048 259398
rect 334448 259954 334768 259986
rect 334448 259718 334490 259954
rect 334726 259718 334768 259954
rect 334448 259634 334768 259718
rect 334448 259398 334490 259634
rect 334726 259398 334768 259634
rect 334448 259366 334768 259398
rect 365168 259954 365488 259986
rect 365168 259718 365210 259954
rect 365446 259718 365488 259954
rect 365168 259634 365488 259718
rect 365168 259398 365210 259634
rect 365446 259398 365488 259634
rect 365168 259366 365488 259398
rect 196208 255454 196528 255486
rect 196208 255218 196250 255454
rect 196486 255218 196528 255454
rect 196208 255134 196528 255218
rect 196208 254898 196250 255134
rect 196486 254898 196528 255134
rect 196208 254866 196528 254898
rect 226928 255454 227248 255486
rect 226928 255218 226970 255454
rect 227206 255218 227248 255454
rect 226928 255134 227248 255218
rect 226928 254898 226970 255134
rect 227206 254898 227248 255134
rect 226928 254866 227248 254898
rect 257648 255454 257968 255486
rect 257648 255218 257690 255454
rect 257926 255218 257968 255454
rect 257648 255134 257968 255218
rect 257648 254898 257690 255134
rect 257926 254898 257968 255134
rect 257648 254866 257968 254898
rect 288368 255454 288688 255486
rect 288368 255218 288410 255454
rect 288646 255218 288688 255454
rect 288368 255134 288688 255218
rect 288368 254898 288410 255134
rect 288646 254898 288688 255134
rect 288368 254866 288688 254898
rect 319088 255454 319408 255486
rect 319088 255218 319130 255454
rect 319366 255218 319408 255454
rect 319088 255134 319408 255218
rect 319088 254898 319130 255134
rect 319366 254898 319408 255134
rect 319088 254866 319408 254898
rect 349808 255454 350128 255486
rect 349808 255218 349850 255454
rect 350086 255218 350128 255454
rect 349808 255134 350128 255218
rect 349808 254898 349850 255134
rect 350086 254898 350128 255134
rect 349808 254866 350128 254898
rect 380528 255454 380848 255486
rect 380528 255218 380570 255454
rect 380806 255218 380848 255454
rect 380528 255134 380848 255218
rect 380528 254898 380570 255134
rect 380806 254898 380848 255134
rect 380528 254866 380848 254898
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 211568 223954 211888 223986
rect 211568 223718 211610 223954
rect 211846 223718 211888 223954
rect 211568 223634 211888 223718
rect 211568 223398 211610 223634
rect 211846 223398 211888 223634
rect 211568 223366 211888 223398
rect 242288 223954 242608 223986
rect 242288 223718 242330 223954
rect 242566 223718 242608 223954
rect 242288 223634 242608 223718
rect 242288 223398 242330 223634
rect 242566 223398 242608 223634
rect 242288 223366 242608 223398
rect 273008 223954 273328 223986
rect 273008 223718 273050 223954
rect 273286 223718 273328 223954
rect 273008 223634 273328 223718
rect 273008 223398 273050 223634
rect 273286 223398 273328 223634
rect 273008 223366 273328 223398
rect 303728 223954 304048 223986
rect 303728 223718 303770 223954
rect 304006 223718 304048 223954
rect 303728 223634 304048 223718
rect 303728 223398 303770 223634
rect 304006 223398 304048 223634
rect 303728 223366 304048 223398
rect 334448 223954 334768 223986
rect 334448 223718 334490 223954
rect 334726 223718 334768 223954
rect 334448 223634 334768 223718
rect 334448 223398 334490 223634
rect 334726 223398 334768 223634
rect 334448 223366 334768 223398
rect 365168 223954 365488 223986
rect 365168 223718 365210 223954
rect 365446 223718 365488 223954
rect 365168 223634 365488 223718
rect 365168 223398 365210 223634
rect 365446 223398 365488 223634
rect 365168 223366 365488 223398
rect 196208 219454 196528 219486
rect 196208 219218 196250 219454
rect 196486 219218 196528 219454
rect 196208 219134 196528 219218
rect 196208 218898 196250 219134
rect 196486 218898 196528 219134
rect 196208 218866 196528 218898
rect 226928 219454 227248 219486
rect 226928 219218 226970 219454
rect 227206 219218 227248 219454
rect 226928 219134 227248 219218
rect 226928 218898 226970 219134
rect 227206 218898 227248 219134
rect 226928 218866 227248 218898
rect 257648 219454 257968 219486
rect 257648 219218 257690 219454
rect 257926 219218 257968 219454
rect 257648 219134 257968 219218
rect 257648 218898 257690 219134
rect 257926 218898 257968 219134
rect 257648 218866 257968 218898
rect 288368 219454 288688 219486
rect 288368 219218 288410 219454
rect 288646 219218 288688 219454
rect 288368 219134 288688 219218
rect 288368 218898 288410 219134
rect 288646 218898 288688 219134
rect 288368 218866 288688 218898
rect 319088 219454 319408 219486
rect 319088 219218 319130 219454
rect 319366 219218 319408 219454
rect 319088 219134 319408 219218
rect 319088 218898 319130 219134
rect 319366 218898 319408 219134
rect 319088 218866 319408 218898
rect 349808 219454 350128 219486
rect 349808 219218 349850 219454
rect 350086 219218 350128 219454
rect 349808 219134 350128 219218
rect 349808 218898 349850 219134
rect 350086 218898 350128 219134
rect 349808 218866 350128 218898
rect 380528 219454 380848 219486
rect 380528 219218 380570 219454
rect 380806 219218 380848 219454
rect 380528 219134 380848 219218
rect 380528 218898 380570 219134
rect 380806 218898 380848 219134
rect 380528 218866 380848 218898
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 211568 187954 211888 187986
rect 211568 187718 211610 187954
rect 211846 187718 211888 187954
rect 211568 187634 211888 187718
rect 211568 187398 211610 187634
rect 211846 187398 211888 187634
rect 211568 187366 211888 187398
rect 242288 187954 242608 187986
rect 242288 187718 242330 187954
rect 242566 187718 242608 187954
rect 242288 187634 242608 187718
rect 242288 187398 242330 187634
rect 242566 187398 242608 187634
rect 242288 187366 242608 187398
rect 273008 187954 273328 187986
rect 273008 187718 273050 187954
rect 273286 187718 273328 187954
rect 273008 187634 273328 187718
rect 273008 187398 273050 187634
rect 273286 187398 273328 187634
rect 273008 187366 273328 187398
rect 303728 187954 304048 187986
rect 303728 187718 303770 187954
rect 304006 187718 304048 187954
rect 303728 187634 304048 187718
rect 303728 187398 303770 187634
rect 304006 187398 304048 187634
rect 303728 187366 304048 187398
rect 334448 187954 334768 187986
rect 334448 187718 334490 187954
rect 334726 187718 334768 187954
rect 334448 187634 334768 187718
rect 334448 187398 334490 187634
rect 334726 187398 334768 187634
rect 334448 187366 334768 187398
rect 365168 187954 365488 187986
rect 365168 187718 365210 187954
rect 365446 187718 365488 187954
rect 365168 187634 365488 187718
rect 365168 187398 365210 187634
rect 365446 187398 365488 187634
rect 365168 187366 365488 187398
rect 196208 183454 196528 183486
rect 196208 183218 196250 183454
rect 196486 183218 196528 183454
rect 196208 183134 196528 183218
rect 196208 182898 196250 183134
rect 196486 182898 196528 183134
rect 196208 182866 196528 182898
rect 226928 183454 227248 183486
rect 226928 183218 226970 183454
rect 227206 183218 227248 183454
rect 226928 183134 227248 183218
rect 226928 182898 226970 183134
rect 227206 182898 227248 183134
rect 226928 182866 227248 182898
rect 257648 183454 257968 183486
rect 257648 183218 257690 183454
rect 257926 183218 257968 183454
rect 257648 183134 257968 183218
rect 257648 182898 257690 183134
rect 257926 182898 257968 183134
rect 257648 182866 257968 182898
rect 288368 183454 288688 183486
rect 288368 183218 288410 183454
rect 288646 183218 288688 183454
rect 288368 183134 288688 183218
rect 288368 182898 288410 183134
rect 288646 182898 288688 183134
rect 288368 182866 288688 182898
rect 319088 183454 319408 183486
rect 319088 183218 319130 183454
rect 319366 183218 319408 183454
rect 319088 183134 319408 183218
rect 319088 182898 319130 183134
rect 319366 182898 319408 183134
rect 319088 182866 319408 182898
rect 349808 183454 350128 183486
rect 349808 183218 349850 183454
rect 350086 183218 350128 183454
rect 349808 183134 350128 183218
rect 349808 182898 349850 183134
rect 350086 182898 350128 183134
rect 349808 182866 350128 182898
rect 380528 183454 380848 183486
rect 380528 183218 380570 183454
rect 380806 183218 380848 183454
rect 380528 183134 380848 183218
rect 380528 182898 380570 183134
rect 380806 182898 380848 183134
rect 380528 182866 380848 182898
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 211568 151954 211888 151986
rect 211568 151718 211610 151954
rect 211846 151718 211888 151954
rect 211568 151634 211888 151718
rect 211568 151398 211610 151634
rect 211846 151398 211888 151634
rect 211568 151366 211888 151398
rect 242288 151954 242608 151986
rect 242288 151718 242330 151954
rect 242566 151718 242608 151954
rect 242288 151634 242608 151718
rect 242288 151398 242330 151634
rect 242566 151398 242608 151634
rect 242288 151366 242608 151398
rect 273008 151954 273328 151986
rect 273008 151718 273050 151954
rect 273286 151718 273328 151954
rect 273008 151634 273328 151718
rect 273008 151398 273050 151634
rect 273286 151398 273328 151634
rect 273008 151366 273328 151398
rect 303728 151954 304048 151986
rect 303728 151718 303770 151954
rect 304006 151718 304048 151954
rect 303728 151634 304048 151718
rect 303728 151398 303770 151634
rect 304006 151398 304048 151634
rect 303728 151366 304048 151398
rect 334448 151954 334768 151986
rect 334448 151718 334490 151954
rect 334726 151718 334768 151954
rect 334448 151634 334768 151718
rect 334448 151398 334490 151634
rect 334726 151398 334768 151634
rect 334448 151366 334768 151398
rect 365168 151954 365488 151986
rect 365168 151718 365210 151954
rect 365446 151718 365488 151954
rect 365168 151634 365488 151718
rect 365168 151398 365210 151634
rect 365446 151398 365488 151634
rect 365168 151366 365488 151398
rect 196208 147454 196528 147486
rect 196208 147218 196250 147454
rect 196486 147218 196528 147454
rect 196208 147134 196528 147218
rect 196208 146898 196250 147134
rect 196486 146898 196528 147134
rect 196208 146866 196528 146898
rect 226928 147454 227248 147486
rect 226928 147218 226970 147454
rect 227206 147218 227248 147454
rect 226928 147134 227248 147218
rect 226928 146898 226970 147134
rect 227206 146898 227248 147134
rect 226928 146866 227248 146898
rect 257648 147454 257968 147486
rect 257648 147218 257690 147454
rect 257926 147218 257968 147454
rect 257648 147134 257968 147218
rect 257648 146898 257690 147134
rect 257926 146898 257968 147134
rect 257648 146866 257968 146898
rect 288368 147454 288688 147486
rect 288368 147218 288410 147454
rect 288646 147218 288688 147454
rect 288368 147134 288688 147218
rect 288368 146898 288410 147134
rect 288646 146898 288688 147134
rect 288368 146866 288688 146898
rect 319088 147454 319408 147486
rect 319088 147218 319130 147454
rect 319366 147218 319408 147454
rect 319088 147134 319408 147218
rect 319088 146898 319130 147134
rect 319366 146898 319408 147134
rect 319088 146866 319408 146898
rect 349808 147454 350128 147486
rect 349808 147218 349850 147454
rect 350086 147218 350128 147454
rect 349808 147134 350128 147218
rect 349808 146898 349850 147134
rect 350086 146898 350128 147134
rect 349808 146866 350128 146898
rect 380528 147454 380848 147486
rect 380528 147218 380570 147454
rect 380806 147218 380848 147454
rect 380528 147134 380848 147218
rect 380528 146898 380570 147134
rect 380806 146898 380848 147134
rect 380528 146866 380848 146898
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 211568 115954 211888 115986
rect 211568 115718 211610 115954
rect 211846 115718 211888 115954
rect 211568 115634 211888 115718
rect 211568 115398 211610 115634
rect 211846 115398 211888 115634
rect 211568 115366 211888 115398
rect 242288 115954 242608 115986
rect 242288 115718 242330 115954
rect 242566 115718 242608 115954
rect 242288 115634 242608 115718
rect 242288 115398 242330 115634
rect 242566 115398 242608 115634
rect 242288 115366 242608 115398
rect 273008 115954 273328 115986
rect 273008 115718 273050 115954
rect 273286 115718 273328 115954
rect 273008 115634 273328 115718
rect 273008 115398 273050 115634
rect 273286 115398 273328 115634
rect 273008 115366 273328 115398
rect 303728 115954 304048 115986
rect 303728 115718 303770 115954
rect 304006 115718 304048 115954
rect 303728 115634 304048 115718
rect 303728 115398 303770 115634
rect 304006 115398 304048 115634
rect 303728 115366 304048 115398
rect 334448 115954 334768 115986
rect 334448 115718 334490 115954
rect 334726 115718 334768 115954
rect 334448 115634 334768 115718
rect 334448 115398 334490 115634
rect 334726 115398 334768 115634
rect 334448 115366 334768 115398
rect 365168 115954 365488 115986
rect 365168 115718 365210 115954
rect 365446 115718 365488 115954
rect 365168 115634 365488 115718
rect 365168 115398 365210 115634
rect 365446 115398 365488 115634
rect 365168 115366 365488 115398
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 84454 191414 108000
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 88954 195914 108000
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 93454 200414 108000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 97954 204914 108000
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 102454 209414 108000
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 106954 213914 108000
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 108000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 79954 222914 108000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 108000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 108000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 108000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 97954 240914 108000
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 102454 245414 108000
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 106954 249914 108000
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 75454 254414 108000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 79954 258914 108000
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 84454 263414 108000
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 88954 267914 108000
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 93454 272414 108000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 97954 276914 108000
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 102454 281414 108000
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 106954 285914 108000
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 75454 290414 108000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 79954 294914 108000
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 84454 299414 108000
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 88954 303914 108000
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 93454 308414 108000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 97954 312914 108000
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 102454 317414 108000
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 106954 321914 108000
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 108000
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 108000
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 84454 335414 108000
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 88954 339914 108000
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 93454 344414 108000
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 97954 348914 108000
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 102454 353414 108000
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 106954 357914 108000
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 75454 362414 108000
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 79954 366914 108000
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 84454 371414 108000
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 88954 375914 108000
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 93454 380414 108000
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 97954 384914 108000
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 102454 389414 108000
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 106954 393914 108000
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 211610 367718 211846 367954
rect 211610 367398 211846 367634
rect 242330 367718 242566 367954
rect 242330 367398 242566 367634
rect 273050 367718 273286 367954
rect 273050 367398 273286 367634
rect 303770 367718 304006 367954
rect 303770 367398 304006 367634
rect 334490 367718 334726 367954
rect 334490 367398 334726 367634
rect 365210 367718 365446 367954
rect 365210 367398 365446 367634
rect 196250 363218 196486 363454
rect 196250 362898 196486 363134
rect 226970 363218 227206 363454
rect 226970 362898 227206 363134
rect 257690 363218 257926 363454
rect 257690 362898 257926 363134
rect 288410 363218 288646 363454
rect 288410 362898 288646 363134
rect 319130 363218 319366 363454
rect 319130 362898 319366 363134
rect 349850 363218 350086 363454
rect 349850 362898 350086 363134
rect 380570 363218 380806 363454
rect 380570 362898 380806 363134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 211610 331718 211846 331954
rect 211610 331398 211846 331634
rect 242330 331718 242566 331954
rect 242330 331398 242566 331634
rect 273050 331718 273286 331954
rect 273050 331398 273286 331634
rect 303770 331718 304006 331954
rect 303770 331398 304006 331634
rect 334490 331718 334726 331954
rect 334490 331398 334726 331634
rect 365210 331718 365446 331954
rect 365210 331398 365446 331634
rect 196250 327218 196486 327454
rect 196250 326898 196486 327134
rect 226970 327218 227206 327454
rect 226970 326898 227206 327134
rect 257690 327218 257926 327454
rect 257690 326898 257926 327134
rect 288410 327218 288646 327454
rect 288410 326898 288646 327134
rect 319130 327218 319366 327454
rect 319130 326898 319366 327134
rect 349850 327218 350086 327454
rect 349850 326898 350086 327134
rect 380570 327218 380806 327454
rect 380570 326898 380806 327134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 211610 295718 211846 295954
rect 211610 295398 211846 295634
rect 242330 295718 242566 295954
rect 242330 295398 242566 295634
rect 273050 295718 273286 295954
rect 273050 295398 273286 295634
rect 303770 295718 304006 295954
rect 303770 295398 304006 295634
rect 334490 295718 334726 295954
rect 334490 295398 334726 295634
rect 365210 295718 365446 295954
rect 365210 295398 365446 295634
rect 196250 291218 196486 291454
rect 196250 290898 196486 291134
rect 226970 291218 227206 291454
rect 226970 290898 227206 291134
rect 257690 291218 257926 291454
rect 257690 290898 257926 291134
rect 288410 291218 288646 291454
rect 288410 290898 288646 291134
rect 319130 291218 319366 291454
rect 319130 290898 319366 291134
rect 349850 291218 350086 291454
rect 349850 290898 350086 291134
rect 380570 291218 380806 291454
rect 380570 290898 380806 291134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 211610 259718 211846 259954
rect 211610 259398 211846 259634
rect 242330 259718 242566 259954
rect 242330 259398 242566 259634
rect 273050 259718 273286 259954
rect 273050 259398 273286 259634
rect 303770 259718 304006 259954
rect 303770 259398 304006 259634
rect 334490 259718 334726 259954
rect 334490 259398 334726 259634
rect 365210 259718 365446 259954
rect 365210 259398 365446 259634
rect 196250 255218 196486 255454
rect 196250 254898 196486 255134
rect 226970 255218 227206 255454
rect 226970 254898 227206 255134
rect 257690 255218 257926 255454
rect 257690 254898 257926 255134
rect 288410 255218 288646 255454
rect 288410 254898 288646 255134
rect 319130 255218 319366 255454
rect 319130 254898 319366 255134
rect 349850 255218 350086 255454
rect 349850 254898 350086 255134
rect 380570 255218 380806 255454
rect 380570 254898 380806 255134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 211610 223718 211846 223954
rect 211610 223398 211846 223634
rect 242330 223718 242566 223954
rect 242330 223398 242566 223634
rect 273050 223718 273286 223954
rect 273050 223398 273286 223634
rect 303770 223718 304006 223954
rect 303770 223398 304006 223634
rect 334490 223718 334726 223954
rect 334490 223398 334726 223634
rect 365210 223718 365446 223954
rect 365210 223398 365446 223634
rect 196250 219218 196486 219454
rect 196250 218898 196486 219134
rect 226970 219218 227206 219454
rect 226970 218898 227206 219134
rect 257690 219218 257926 219454
rect 257690 218898 257926 219134
rect 288410 219218 288646 219454
rect 288410 218898 288646 219134
rect 319130 219218 319366 219454
rect 319130 218898 319366 219134
rect 349850 219218 350086 219454
rect 349850 218898 350086 219134
rect 380570 219218 380806 219454
rect 380570 218898 380806 219134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 211610 187718 211846 187954
rect 211610 187398 211846 187634
rect 242330 187718 242566 187954
rect 242330 187398 242566 187634
rect 273050 187718 273286 187954
rect 273050 187398 273286 187634
rect 303770 187718 304006 187954
rect 303770 187398 304006 187634
rect 334490 187718 334726 187954
rect 334490 187398 334726 187634
rect 365210 187718 365446 187954
rect 365210 187398 365446 187634
rect 196250 183218 196486 183454
rect 196250 182898 196486 183134
rect 226970 183218 227206 183454
rect 226970 182898 227206 183134
rect 257690 183218 257926 183454
rect 257690 182898 257926 183134
rect 288410 183218 288646 183454
rect 288410 182898 288646 183134
rect 319130 183218 319366 183454
rect 319130 182898 319366 183134
rect 349850 183218 350086 183454
rect 349850 182898 350086 183134
rect 380570 183218 380806 183454
rect 380570 182898 380806 183134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 211610 151718 211846 151954
rect 211610 151398 211846 151634
rect 242330 151718 242566 151954
rect 242330 151398 242566 151634
rect 273050 151718 273286 151954
rect 273050 151398 273286 151634
rect 303770 151718 304006 151954
rect 303770 151398 304006 151634
rect 334490 151718 334726 151954
rect 334490 151398 334726 151634
rect 365210 151718 365446 151954
rect 365210 151398 365446 151634
rect 196250 147218 196486 147454
rect 196250 146898 196486 147134
rect 226970 147218 227206 147454
rect 226970 146898 227206 147134
rect 257690 147218 257926 147454
rect 257690 146898 257926 147134
rect 288410 147218 288646 147454
rect 288410 146898 288646 147134
rect 319130 147218 319366 147454
rect 319130 146898 319366 147134
rect 349850 147218 350086 147454
rect 349850 146898 350086 147134
rect 380570 147218 380806 147454
rect 380570 146898 380806 147134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 211610 115718 211846 115954
rect 211610 115398 211846 115634
rect 242330 115718 242566 115954
rect 242330 115398 242566 115634
rect 273050 115718 273286 115954
rect 273050 115398 273286 115634
rect 303770 115718 304006 115954
rect 303770 115398 304006 115634
rect 334490 115718 334726 115954
rect 334490 115398 334726 115634
rect 365210 115718 365446 115954
rect 365210 115398 365446 115634
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 211610 367954
rect 211846 367718 242330 367954
rect 242566 367718 273050 367954
rect 273286 367718 303770 367954
rect 304006 367718 334490 367954
rect 334726 367718 365210 367954
rect 365446 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 211610 367634
rect 211846 367398 242330 367634
rect 242566 367398 273050 367634
rect 273286 367398 303770 367634
rect 304006 367398 334490 367634
rect 334726 367398 365210 367634
rect 365446 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 196250 363454
rect 196486 363218 226970 363454
rect 227206 363218 257690 363454
rect 257926 363218 288410 363454
rect 288646 363218 319130 363454
rect 319366 363218 349850 363454
rect 350086 363218 380570 363454
rect 380806 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 196250 363134
rect 196486 362898 226970 363134
rect 227206 362898 257690 363134
rect 257926 362898 288410 363134
rect 288646 362898 319130 363134
rect 319366 362898 349850 363134
rect 350086 362898 380570 363134
rect 380806 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 211610 331954
rect 211846 331718 242330 331954
rect 242566 331718 273050 331954
rect 273286 331718 303770 331954
rect 304006 331718 334490 331954
rect 334726 331718 365210 331954
rect 365446 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 211610 331634
rect 211846 331398 242330 331634
rect 242566 331398 273050 331634
rect 273286 331398 303770 331634
rect 304006 331398 334490 331634
rect 334726 331398 365210 331634
rect 365446 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 196250 327454
rect 196486 327218 226970 327454
rect 227206 327218 257690 327454
rect 257926 327218 288410 327454
rect 288646 327218 319130 327454
rect 319366 327218 349850 327454
rect 350086 327218 380570 327454
rect 380806 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 196250 327134
rect 196486 326898 226970 327134
rect 227206 326898 257690 327134
rect 257926 326898 288410 327134
rect 288646 326898 319130 327134
rect 319366 326898 349850 327134
rect 350086 326898 380570 327134
rect 380806 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 211610 295954
rect 211846 295718 242330 295954
rect 242566 295718 273050 295954
rect 273286 295718 303770 295954
rect 304006 295718 334490 295954
rect 334726 295718 365210 295954
rect 365446 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 211610 295634
rect 211846 295398 242330 295634
rect 242566 295398 273050 295634
rect 273286 295398 303770 295634
rect 304006 295398 334490 295634
rect 334726 295398 365210 295634
rect 365446 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 196250 291454
rect 196486 291218 226970 291454
rect 227206 291218 257690 291454
rect 257926 291218 288410 291454
rect 288646 291218 319130 291454
rect 319366 291218 349850 291454
rect 350086 291218 380570 291454
rect 380806 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 196250 291134
rect 196486 290898 226970 291134
rect 227206 290898 257690 291134
rect 257926 290898 288410 291134
rect 288646 290898 319130 291134
rect 319366 290898 349850 291134
rect 350086 290898 380570 291134
rect 380806 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 211610 259954
rect 211846 259718 242330 259954
rect 242566 259718 273050 259954
rect 273286 259718 303770 259954
rect 304006 259718 334490 259954
rect 334726 259718 365210 259954
rect 365446 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 211610 259634
rect 211846 259398 242330 259634
rect 242566 259398 273050 259634
rect 273286 259398 303770 259634
rect 304006 259398 334490 259634
rect 334726 259398 365210 259634
rect 365446 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 196250 255454
rect 196486 255218 226970 255454
rect 227206 255218 257690 255454
rect 257926 255218 288410 255454
rect 288646 255218 319130 255454
rect 319366 255218 349850 255454
rect 350086 255218 380570 255454
rect 380806 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 196250 255134
rect 196486 254898 226970 255134
rect 227206 254898 257690 255134
rect 257926 254898 288410 255134
rect 288646 254898 319130 255134
rect 319366 254898 349850 255134
rect 350086 254898 380570 255134
rect 380806 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 211610 223954
rect 211846 223718 242330 223954
rect 242566 223718 273050 223954
rect 273286 223718 303770 223954
rect 304006 223718 334490 223954
rect 334726 223718 365210 223954
rect 365446 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 211610 223634
rect 211846 223398 242330 223634
rect 242566 223398 273050 223634
rect 273286 223398 303770 223634
rect 304006 223398 334490 223634
rect 334726 223398 365210 223634
rect 365446 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 196250 219454
rect 196486 219218 226970 219454
rect 227206 219218 257690 219454
rect 257926 219218 288410 219454
rect 288646 219218 319130 219454
rect 319366 219218 349850 219454
rect 350086 219218 380570 219454
rect 380806 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 196250 219134
rect 196486 218898 226970 219134
rect 227206 218898 257690 219134
rect 257926 218898 288410 219134
rect 288646 218898 319130 219134
rect 319366 218898 349850 219134
rect 350086 218898 380570 219134
rect 380806 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 211610 187954
rect 211846 187718 242330 187954
rect 242566 187718 273050 187954
rect 273286 187718 303770 187954
rect 304006 187718 334490 187954
rect 334726 187718 365210 187954
rect 365446 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 211610 187634
rect 211846 187398 242330 187634
rect 242566 187398 273050 187634
rect 273286 187398 303770 187634
rect 304006 187398 334490 187634
rect 334726 187398 365210 187634
rect 365446 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 196250 183454
rect 196486 183218 226970 183454
rect 227206 183218 257690 183454
rect 257926 183218 288410 183454
rect 288646 183218 319130 183454
rect 319366 183218 349850 183454
rect 350086 183218 380570 183454
rect 380806 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 196250 183134
rect 196486 182898 226970 183134
rect 227206 182898 257690 183134
rect 257926 182898 288410 183134
rect 288646 182898 319130 183134
rect 319366 182898 349850 183134
rect 350086 182898 380570 183134
rect 380806 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 211610 151954
rect 211846 151718 242330 151954
rect 242566 151718 273050 151954
rect 273286 151718 303770 151954
rect 304006 151718 334490 151954
rect 334726 151718 365210 151954
rect 365446 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 211610 151634
rect 211846 151398 242330 151634
rect 242566 151398 273050 151634
rect 273286 151398 303770 151634
rect 304006 151398 334490 151634
rect 334726 151398 365210 151634
rect 365446 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 196250 147454
rect 196486 147218 226970 147454
rect 227206 147218 257690 147454
rect 257926 147218 288410 147454
rect 288646 147218 319130 147454
rect 319366 147218 349850 147454
rect 350086 147218 380570 147454
rect 380806 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 196250 147134
rect 196486 146898 226970 147134
rect 227206 146898 257690 147134
rect 257926 146898 288410 147134
rect 288646 146898 319130 147134
rect 319366 146898 349850 147134
rect 350086 146898 380570 147134
rect 380806 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 211610 115954
rect 211846 115718 242330 115954
rect 242566 115718 273050 115954
rect 273286 115718 303770 115954
rect 304006 115718 334490 115954
rect 334726 115718 365210 115954
rect 365446 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 211610 115634
rect 211846 115398 242330 115634
rect 242566 115398 273050 115634
rect 273286 115398 303770 115634
rect 304006 115398 334490 115634
rect 334726 115398 365210 115634
rect 365446 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 192000 0 1 110000
box 0 0 200000 280000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 108000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 392000 218414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 108000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 392000 254414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 108000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 392000 290414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 108000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 392000 326414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 108000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 392000 362414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 392000 191414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 392000 227414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 392000 263414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 392000 299414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 392000 335414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 108000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 392000 371414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 392000 200414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 392000 236414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 392000 272414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 392000 308414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 392000 344414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 108000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 392000 380414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 392000 209414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 392000 245414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 392000 281414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 392000 317414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 392000 353414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 108000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 392000 389414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 392000 204914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 392000 240914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 392000 276914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 392000 312914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 392000 348914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 108000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 392000 384914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 392000 213914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 392000 249914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 392000 285914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 392000 321914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 392000 357914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 108000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 392000 393914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 108000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 392000 222914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 108000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 392000 258914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 108000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 392000 294914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 108000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 392000 330914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 108000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 392000 366914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 392000 195914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 392000 231914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 392000 267914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 392000 303914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 392000 339914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 108000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 392000 375914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
