magic
tech sky130A
magscale 1 2
timestamp 1654529215
<< obsli1 >>
rect 1104 2159 198812 277457
<< obsm1 >>
rect 198 1436 199810 277488
<< metal2 >>
rect 3698 279200 3754 280000
rect 11058 279200 11114 280000
rect 18510 279200 18566 280000
rect 25870 279200 25926 280000
rect 33322 279200 33378 280000
rect 40682 279200 40738 280000
rect 48134 279200 48190 280000
rect 55494 279200 55550 280000
rect 62946 279200 63002 280000
rect 70306 279200 70362 280000
rect 77758 279200 77814 280000
rect 85118 279200 85174 280000
rect 92570 279200 92626 280000
rect 99930 279200 99986 280000
rect 107382 279200 107438 280000
rect 114742 279200 114798 280000
rect 122194 279200 122250 280000
rect 129554 279200 129610 280000
rect 137006 279200 137062 280000
rect 144366 279200 144422 280000
rect 151818 279200 151874 280000
rect 159178 279200 159234 280000
rect 166630 279200 166686 280000
rect 173990 279200 174046 280000
rect 181442 279200 181498 280000
rect 188802 279200 188858 280000
rect 196254 279200 196310 280000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61842 0 61898 800
rect 62210 0 62266 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89810 0 89866 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91466 0 91522 800
rect 91834 0 91890 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103978 0 104034 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109314 0 109370 800
rect 109682 0 109738 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 119066 0 119122 800
rect 119434 0 119490 800
rect 119802 0 119858 800
rect 120262 0 120318 800
rect 120630 0 120686 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126702 0 126758 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148598 0 148654 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157522 0 157578 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161662 0 161718 800
rect 162030 0 162086 800
rect 162398 0 162454 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164882 0 164938 800
rect 165250 0 165306 800
rect 165710 0 165766 800
rect 166078 0 166134 800
rect 166446 0 166502 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167734 0 167790 800
rect 168102 0 168158 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169758 0 169814 800
rect 170126 0 170182 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172610 0 172666 800
rect 172978 0 173034 800
rect 173346 0 173402 800
rect 173806 0 173862 800
rect 174174 0 174230 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176658 0 176714 800
rect 177026 0 177082 800
rect 177486 0 177542 800
rect 177854 0 177910 800
rect 178222 0 178278 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179510 0 179566 800
rect 179878 0 179934 800
rect 180246 0 180302 800
rect 180706 0 180762 800
rect 181074 0 181130 800
rect 181534 0 181590 800
rect 181902 0 181958 800
rect 182270 0 182326 800
rect 182730 0 182786 800
rect 183098 0 183154 800
rect 183558 0 183614 800
rect 183926 0 183982 800
rect 184386 0 184442 800
rect 184754 0 184810 800
rect 185122 0 185178 800
rect 185582 0 185638 800
rect 185950 0 186006 800
rect 186410 0 186466 800
rect 186778 0 186834 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 187974 0 188030 800
rect 188434 0 188490 800
rect 188802 0 188858 800
rect 189170 0 189226 800
rect 189630 0 189686 800
rect 189998 0 190054 800
rect 190458 0 190514 800
rect 190826 0 190882 800
rect 191194 0 191250 800
rect 191654 0 191710 800
rect 192022 0 192078 800
rect 192482 0 192538 800
rect 192850 0 192906 800
rect 193310 0 193366 800
rect 193678 0 193734 800
rect 194046 0 194102 800
rect 194506 0 194562 800
rect 194874 0 194930 800
rect 195334 0 195390 800
rect 195702 0 195758 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197726 0 197782 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199750 0 199806 800
<< obsm2 >>
rect 204 279144 3642 279200
rect 3810 279144 11002 279200
rect 11170 279144 18454 279200
rect 18622 279144 25814 279200
rect 25982 279144 33266 279200
rect 33434 279144 40626 279200
rect 40794 279144 48078 279200
rect 48246 279144 55438 279200
rect 55606 279144 62890 279200
rect 63058 279144 70250 279200
rect 70418 279144 77702 279200
rect 77870 279144 85062 279200
rect 85230 279144 92514 279200
rect 92682 279144 99874 279200
rect 100042 279144 107326 279200
rect 107494 279144 114686 279200
rect 114854 279144 122138 279200
rect 122306 279144 129498 279200
rect 129666 279144 136950 279200
rect 137118 279144 144310 279200
rect 144478 279144 151762 279200
rect 151930 279144 159122 279200
rect 159290 279144 166574 279200
rect 166742 279144 173934 279200
rect 174102 279144 181386 279200
rect 181554 279144 188746 279200
rect 188914 279144 196198 279200
rect 196366 279144 199804 279200
rect 204 856 199804 279144
rect 314 734 514 856
rect 682 734 882 856
rect 1050 734 1342 856
rect 1510 734 1710 856
rect 1878 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3366 856
rect 3534 734 3734 856
rect 3902 734 4194 856
rect 4362 734 4562 856
rect 4730 734 4930 856
rect 5098 734 5390 856
rect 5558 734 5758 856
rect 5926 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7414 856
rect 7582 734 7782 856
rect 7950 734 8242 856
rect 8410 734 8610 856
rect 8778 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9806 856
rect 9974 734 10266 856
rect 10434 734 10634 856
rect 10802 734 11094 856
rect 11262 734 11462 856
rect 11630 734 11830 856
rect 11998 734 12290 856
rect 12458 734 12658 856
rect 12826 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14314 856
rect 14482 734 14682 856
rect 14850 734 15142 856
rect 15310 734 15510 856
rect 15678 734 15878 856
rect 16046 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17166 856
rect 17334 734 17534 856
rect 17702 734 17994 856
rect 18162 734 18362 856
rect 18530 734 18730 856
rect 18898 734 19190 856
rect 19358 734 19558 856
rect 19726 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20754 856
rect 20922 734 21214 856
rect 21382 734 21582 856
rect 21750 734 22042 856
rect 22210 734 22410 856
rect 22578 734 22778 856
rect 22946 734 23238 856
rect 23406 734 23606 856
rect 23774 734 24066 856
rect 24234 734 24434 856
rect 24602 734 24802 856
rect 24970 734 25262 856
rect 25430 734 25630 856
rect 25798 734 26090 856
rect 26258 734 26458 856
rect 26626 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27654 856
rect 27822 734 28114 856
rect 28282 734 28482 856
rect 28650 734 28942 856
rect 29110 734 29310 856
rect 29478 734 29678 856
rect 29846 734 30138 856
rect 30306 734 30506 856
rect 30674 734 30966 856
rect 31134 734 31334 856
rect 31502 734 31702 856
rect 31870 734 32162 856
rect 32330 734 32530 856
rect 32698 734 32990 856
rect 33158 734 33358 856
rect 33526 734 33818 856
rect 33986 734 34186 856
rect 34354 734 34554 856
rect 34722 734 35014 856
rect 35182 734 35382 856
rect 35550 734 35842 856
rect 36010 734 36210 856
rect 36378 734 36578 856
rect 36746 734 37038 856
rect 37206 734 37406 856
rect 37574 734 37866 856
rect 38034 734 38234 856
rect 38402 734 38602 856
rect 38770 734 39062 856
rect 39230 734 39430 856
rect 39598 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40626 856
rect 40794 734 41086 856
rect 41254 734 41454 856
rect 41622 734 41914 856
rect 42082 734 42282 856
rect 42450 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43478 856
rect 43646 734 43938 856
rect 44106 734 44306 856
rect 44474 734 44766 856
rect 44934 734 45134 856
rect 45302 734 45502 856
rect 45670 734 45962 856
rect 46130 734 46330 856
rect 46498 734 46790 856
rect 46958 734 47158 856
rect 47326 734 47526 856
rect 47694 734 47986 856
rect 48154 734 48354 856
rect 48522 734 48814 856
rect 48982 734 49182 856
rect 49350 734 49550 856
rect 49718 734 50010 856
rect 50178 734 50378 856
rect 50546 734 50838 856
rect 51006 734 51206 856
rect 51374 734 51666 856
rect 51834 734 52034 856
rect 52202 734 52402 856
rect 52570 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53690 856
rect 53858 734 54058 856
rect 54226 734 54426 856
rect 54594 734 54886 856
rect 55054 734 55254 856
rect 55422 734 55714 856
rect 55882 734 56082 856
rect 56250 734 56450 856
rect 56618 734 56910 856
rect 57078 734 57278 856
rect 57446 734 57738 856
rect 57906 734 58106 856
rect 58274 734 58566 856
rect 58734 734 58934 856
rect 59102 734 59302 856
rect 59470 734 59762 856
rect 59930 734 60130 856
rect 60298 734 60590 856
rect 60758 734 60958 856
rect 61126 734 61326 856
rect 61494 734 61786 856
rect 61954 734 62154 856
rect 62322 734 62614 856
rect 62782 734 62982 856
rect 63150 734 63350 856
rect 63518 734 63810 856
rect 63978 734 64178 856
rect 64346 734 64638 856
rect 64806 734 65006 856
rect 65174 734 65374 856
rect 65542 734 65834 856
rect 66002 734 66202 856
rect 66370 734 66662 856
rect 66830 734 67030 856
rect 67198 734 67490 856
rect 67658 734 67858 856
rect 68026 734 68226 856
rect 68394 734 68686 856
rect 68854 734 69054 856
rect 69222 734 69514 856
rect 69682 734 69882 856
rect 70050 734 70250 856
rect 70418 734 70710 856
rect 70878 734 71078 856
rect 71246 734 71538 856
rect 71706 734 71906 856
rect 72074 734 72274 856
rect 72442 734 72734 856
rect 72902 734 73102 856
rect 73270 734 73562 856
rect 73730 734 73930 856
rect 74098 734 74298 856
rect 74466 734 74758 856
rect 74926 734 75126 856
rect 75294 734 75586 856
rect 75754 734 75954 856
rect 76122 734 76414 856
rect 76582 734 76782 856
rect 76950 734 77150 856
rect 77318 734 77610 856
rect 77778 734 77978 856
rect 78146 734 78438 856
rect 78606 734 78806 856
rect 78974 734 79174 856
rect 79342 734 79634 856
rect 79802 734 80002 856
rect 80170 734 80462 856
rect 80630 734 80830 856
rect 80998 734 81198 856
rect 81366 734 81658 856
rect 81826 734 82026 856
rect 82194 734 82486 856
rect 82654 734 82854 856
rect 83022 734 83222 856
rect 83390 734 83682 856
rect 83850 734 84050 856
rect 84218 734 84510 856
rect 84678 734 84878 856
rect 85046 734 85338 856
rect 85506 734 85706 856
rect 85874 734 86074 856
rect 86242 734 86534 856
rect 86702 734 86902 856
rect 87070 734 87362 856
rect 87530 734 87730 856
rect 87898 734 88098 856
rect 88266 734 88558 856
rect 88726 734 88926 856
rect 89094 734 89386 856
rect 89554 734 89754 856
rect 89922 734 90122 856
rect 90290 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91410 856
rect 91578 734 91778 856
rect 91946 734 92238 856
rect 92406 734 92606 856
rect 92774 734 92974 856
rect 93142 734 93434 856
rect 93602 734 93802 856
rect 93970 734 94262 856
rect 94430 734 94630 856
rect 94798 734 94998 856
rect 95166 734 95458 856
rect 95626 734 95826 856
rect 95994 734 96286 856
rect 96454 734 96654 856
rect 96822 734 97022 856
rect 97190 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98310 856
rect 98478 734 98678 856
rect 98846 734 99046 856
rect 99214 734 99506 856
rect 99674 734 99874 856
rect 100042 734 100334 856
rect 100502 734 100702 856
rect 100870 734 101162 856
rect 101330 734 101530 856
rect 101698 734 101898 856
rect 102066 734 102358 856
rect 102526 734 102726 856
rect 102894 734 103186 856
rect 103354 734 103554 856
rect 103722 734 103922 856
rect 104090 734 104382 856
rect 104550 734 104750 856
rect 104918 734 105210 856
rect 105378 734 105578 856
rect 105746 734 105946 856
rect 106114 734 106406 856
rect 106574 734 106774 856
rect 106942 734 107234 856
rect 107402 734 107602 856
rect 107770 734 107970 856
rect 108138 734 108430 856
rect 108598 734 108798 856
rect 108966 734 109258 856
rect 109426 734 109626 856
rect 109794 734 110086 856
rect 110254 734 110454 856
rect 110622 734 110822 856
rect 110990 734 111282 856
rect 111450 734 111650 856
rect 111818 734 112110 856
rect 112278 734 112478 856
rect 112646 734 112846 856
rect 113014 734 113306 856
rect 113474 734 113674 856
rect 113842 734 114134 856
rect 114302 734 114502 856
rect 114670 734 114870 856
rect 115038 734 115330 856
rect 115498 734 115698 856
rect 115866 734 116158 856
rect 116326 734 116526 856
rect 116694 734 116986 856
rect 117154 734 117354 856
rect 117522 734 117722 856
rect 117890 734 118182 856
rect 118350 734 118550 856
rect 118718 734 119010 856
rect 119178 734 119378 856
rect 119546 734 119746 856
rect 119914 734 120206 856
rect 120374 734 120574 856
rect 120742 734 121034 856
rect 121202 734 121402 856
rect 121570 734 121770 856
rect 121938 734 122230 856
rect 122398 734 122598 856
rect 122766 734 123058 856
rect 123226 734 123426 856
rect 123594 734 123794 856
rect 123962 734 124254 856
rect 124422 734 124622 856
rect 124790 734 125082 856
rect 125250 734 125450 856
rect 125618 734 125910 856
rect 126078 734 126278 856
rect 126446 734 126646 856
rect 126814 734 127106 856
rect 127274 734 127474 856
rect 127642 734 127934 856
rect 128102 734 128302 856
rect 128470 734 128670 856
rect 128838 734 129130 856
rect 129298 734 129498 856
rect 129666 734 129958 856
rect 130126 734 130326 856
rect 130494 734 130694 856
rect 130862 734 131154 856
rect 131322 734 131522 856
rect 131690 734 131982 856
rect 132150 734 132350 856
rect 132518 734 132718 856
rect 132886 734 133178 856
rect 133346 734 133546 856
rect 133714 734 134006 856
rect 134174 734 134374 856
rect 134542 734 134834 856
rect 135002 734 135202 856
rect 135370 734 135570 856
rect 135738 734 136030 856
rect 136198 734 136398 856
rect 136566 734 136858 856
rect 137026 734 137226 856
rect 137394 734 137594 856
rect 137762 734 138054 856
rect 138222 734 138422 856
rect 138590 734 138882 856
rect 139050 734 139250 856
rect 139418 734 139618 856
rect 139786 734 140078 856
rect 140246 734 140446 856
rect 140614 734 140906 856
rect 141074 734 141274 856
rect 141442 734 141642 856
rect 141810 734 142102 856
rect 142270 734 142470 856
rect 142638 734 142930 856
rect 143098 734 143298 856
rect 143466 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144494 856
rect 144662 734 144954 856
rect 145122 734 145322 856
rect 145490 734 145782 856
rect 145950 734 146150 856
rect 146318 734 146518 856
rect 146686 734 146978 856
rect 147146 734 147346 856
rect 147514 734 147806 856
rect 147974 734 148174 856
rect 148342 734 148542 856
rect 148710 734 149002 856
rect 149170 734 149370 856
rect 149538 734 149830 856
rect 149998 734 150198 856
rect 150366 734 150658 856
rect 150826 734 151026 856
rect 151194 734 151394 856
rect 151562 734 151854 856
rect 152022 734 152222 856
rect 152390 734 152682 856
rect 152850 734 153050 856
rect 153218 734 153418 856
rect 153586 734 153878 856
rect 154046 734 154246 856
rect 154414 734 154706 856
rect 154874 734 155074 856
rect 155242 734 155442 856
rect 155610 734 155902 856
rect 156070 734 156270 856
rect 156438 734 156730 856
rect 156898 734 157098 856
rect 157266 734 157466 856
rect 157634 734 157926 856
rect 158094 734 158294 856
rect 158462 734 158754 856
rect 158922 734 159122 856
rect 159290 734 159582 856
rect 159750 734 159950 856
rect 160118 734 160318 856
rect 160486 734 160778 856
rect 160946 734 161146 856
rect 161314 734 161606 856
rect 161774 734 161974 856
rect 162142 734 162342 856
rect 162510 734 162802 856
rect 162970 734 163170 856
rect 163338 734 163630 856
rect 163798 734 163998 856
rect 164166 734 164366 856
rect 164534 734 164826 856
rect 164994 734 165194 856
rect 165362 734 165654 856
rect 165822 734 166022 856
rect 166190 734 166390 856
rect 166558 734 166850 856
rect 167018 734 167218 856
rect 167386 734 167678 856
rect 167846 734 168046 856
rect 168214 734 168506 856
rect 168674 734 168874 856
rect 169042 734 169242 856
rect 169410 734 169702 856
rect 169870 734 170070 856
rect 170238 734 170530 856
rect 170698 734 170898 856
rect 171066 734 171266 856
rect 171434 734 171726 856
rect 171894 734 172094 856
rect 172262 734 172554 856
rect 172722 734 172922 856
rect 173090 734 173290 856
rect 173458 734 173750 856
rect 173918 734 174118 856
rect 174286 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175406 856
rect 175574 734 175774 856
rect 175942 734 176142 856
rect 176310 734 176602 856
rect 176770 734 176970 856
rect 177138 734 177430 856
rect 177598 734 177798 856
rect 177966 734 178166 856
rect 178334 734 178626 856
rect 178794 734 178994 856
rect 179162 734 179454 856
rect 179622 734 179822 856
rect 179990 734 180190 856
rect 180358 734 180650 856
rect 180818 734 181018 856
rect 181186 734 181478 856
rect 181646 734 181846 856
rect 182014 734 182214 856
rect 182382 734 182674 856
rect 182842 734 183042 856
rect 183210 734 183502 856
rect 183670 734 183870 856
rect 184038 734 184330 856
rect 184498 734 184698 856
rect 184866 734 185066 856
rect 185234 734 185526 856
rect 185694 734 185894 856
rect 186062 734 186354 856
rect 186522 734 186722 856
rect 186890 734 187090 856
rect 187258 734 187550 856
rect 187718 734 187918 856
rect 188086 734 188378 856
rect 188546 734 188746 856
rect 188914 734 189114 856
rect 189282 734 189574 856
rect 189742 734 189942 856
rect 190110 734 190402 856
rect 190570 734 190770 856
rect 190938 734 191138 856
rect 191306 734 191598 856
rect 191766 734 191966 856
rect 192134 734 192426 856
rect 192594 734 192794 856
rect 192962 734 193254 856
rect 193422 734 193622 856
rect 193790 734 193990 856
rect 194158 734 194450 856
rect 194618 734 194818 856
rect 194986 734 195278 856
rect 195446 734 195646 856
rect 195814 734 196014 856
rect 196182 734 196474 856
rect 196642 734 196842 856
rect 197010 734 197302 856
rect 197470 734 197670 856
rect 197838 734 198038 856
rect 198206 734 198498 856
rect 198666 734 198866 856
rect 199034 734 199326 856
rect 199494 734 199694 856
<< metal3 >>
rect 199200 276768 200000 276888
rect 0 276496 800 276616
rect 199200 270512 200000 270632
rect 0 269832 800 269952
rect 199200 264256 200000 264376
rect 0 263168 800 263288
rect 199200 258000 200000 258120
rect 0 256504 800 256624
rect 199200 251880 200000 252000
rect 0 249840 800 249960
rect 199200 245624 200000 245744
rect 0 243176 800 243296
rect 199200 239368 200000 239488
rect 0 236512 800 236632
rect 199200 233112 200000 233232
rect 0 229848 800 229968
rect 199200 226992 200000 227112
rect 0 223184 800 223304
rect 199200 220736 200000 220856
rect 0 216520 800 216640
rect 199200 214480 200000 214600
rect 0 209856 800 209976
rect 199200 208224 200000 208344
rect 0 203192 800 203312
rect 199200 202104 200000 202224
rect 0 196528 800 196648
rect 199200 195848 200000 195968
rect 0 189864 800 189984
rect 199200 189592 200000 189712
rect 0 183200 800 183320
rect 199200 183336 200000 183456
rect 199200 177216 200000 177336
rect 0 176536 800 176656
rect 199200 170960 200000 171080
rect 0 169872 800 169992
rect 199200 164704 200000 164824
rect 0 163208 800 163328
rect 199200 158448 200000 158568
rect 0 156544 800 156664
rect 199200 152328 200000 152448
rect 0 149880 800 150000
rect 199200 146072 200000 146192
rect 0 143216 800 143336
rect 199200 139816 200000 139936
rect 0 136552 800 136672
rect 199200 133560 200000 133680
rect 0 129888 800 130008
rect 199200 127440 200000 127560
rect 0 123224 800 123344
rect 199200 121184 200000 121304
rect 0 116560 800 116680
rect 199200 114928 200000 115048
rect 0 109896 800 110016
rect 199200 108672 200000 108792
rect 0 103232 800 103352
rect 199200 102552 200000 102672
rect 0 96568 800 96688
rect 199200 96296 200000 96416
rect 0 89904 800 90024
rect 199200 90040 200000 90160
rect 199200 83784 200000 83904
rect 0 83240 800 83360
rect 199200 77664 200000 77784
rect 0 76576 800 76696
rect 199200 71408 200000 71528
rect 0 69912 800 70032
rect 199200 65152 200000 65272
rect 0 63248 800 63368
rect 199200 58896 200000 59016
rect 0 56584 800 56704
rect 199200 52776 200000 52896
rect 0 49920 800 50040
rect 199200 46520 200000 46640
rect 0 43256 800 43376
rect 199200 40264 200000 40384
rect 0 36592 800 36712
rect 199200 34008 200000 34128
rect 0 29928 800 30048
rect 199200 27888 200000 28008
rect 0 23264 800 23384
rect 199200 21632 200000 21752
rect 0 16600 800 16720
rect 199200 15376 200000 15496
rect 0 9936 800 10056
rect 199200 9120 200000 9240
rect 0 3272 800 3392
rect 199200 3000 200000 3120
<< obsm3 >>
rect 800 276968 199200 277473
rect 800 276696 199120 276968
rect 880 276688 199120 276696
rect 880 276416 199200 276688
rect 800 270712 199200 276416
rect 800 270432 199120 270712
rect 800 270032 199200 270432
rect 880 269752 199200 270032
rect 800 264456 199200 269752
rect 800 264176 199120 264456
rect 800 263368 199200 264176
rect 880 263088 199200 263368
rect 800 258200 199200 263088
rect 800 257920 199120 258200
rect 800 256704 199200 257920
rect 880 256424 199200 256704
rect 800 252080 199200 256424
rect 800 251800 199120 252080
rect 800 250040 199200 251800
rect 880 249760 199200 250040
rect 800 245824 199200 249760
rect 800 245544 199120 245824
rect 800 243376 199200 245544
rect 880 243096 199200 243376
rect 800 239568 199200 243096
rect 800 239288 199120 239568
rect 800 236712 199200 239288
rect 880 236432 199200 236712
rect 800 233312 199200 236432
rect 800 233032 199120 233312
rect 800 230048 199200 233032
rect 880 229768 199200 230048
rect 800 227192 199200 229768
rect 800 226912 199120 227192
rect 800 223384 199200 226912
rect 880 223104 199200 223384
rect 800 220936 199200 223104
rect 800 220656 199120 220936
rect 800 216720 199200 220656
rect 880 216440 199200 216720
rect 800 214680 199200 216440
rect 800 214400 199120 214680
rect 800 210056 199200 214400
rect 880 209776 199200 210056
rect 800 208424 199200 209776
rect 800 208144 199120 208424
rect 800 203392 199200 208144
rect 880 203112 199200 203392
rect 800 202304 199200 203112
rect 800 202024 199120 202304
rect 800 196728 199200 202024
rect 880 196448 199200 196728
rect 800 196048 199200 196448
rect 800 195768 199120 196048
rect 800 190064 199200 195768
rect 880 189792 199200 190064
rect 880 189784 199120 189792
rect 800 189512 199120 189784
rect 800 183536 199200 189512
rect 800 183400 199120 183536
rect 880 183256 199120 183400
rect 880 183120 199200 183256
rect 800 177416 199200 183120
rect 800 177136 199120 177416
rect 800 176736 199200 177136
rect 880 176456 199200 176736
rect 800 171160 199200 176456
rect 800 170880 199120 171160
rect 800 170072 199200 170880
rect 880 169792 199200 170072
rect 800 164904 199200 169792
rect 800 164624 199120 164904
rect 800 163408 199200 164624
rect 880 163128 199200 163408
rect 800 158648 199200 163128
rect 800 158368 199120 158648
rect 800 156744 199200 158368
rect 880 156464 199200 156744
rect 800 152528 199200 156464
rect 800 152248 199120 152528
rect 800 150080 199200 152248
rect 880 149800 199200 150080
rect 800 146272 199200 149800
rect 800 145992 199120 146272
rect 800 143416 199200 145992
rect 880 143136 199200 143416
rect 800 140016 199200 143136
rect 800 139736 199120 140016
rect 800 136752 199200 139736
rect 880 136472 199200 136752
rect 800 133760 199200 136472
rect 800 133480 199120 133760
rect 800 130088 199200 133480
rect 880 129808 199200 130088
rect 800 127640 199200 129808
rect 800 127360 199120 127640
rect 800 123424 199200 127360
rect 880 123144 199200 123424
rect 800 121384 199200 123144
rect 800 121104 199120 121384
rect 800 116760 199200 121104
rect 880 116480 199200 116760
rect 800 115128 199200 116480
rect 800 114848 199120 115128
rect 800 110096 199200 114848
rect 880 109816 199200 110096
rect 800 108872 199200 109816
rect 800 108592 199120 108872
rect 800 103432 199200 108592
rect 880 103152 199200 103432
rect 800 102752 199200 103152
rect 800 102472 199120 102752
rect 800 96768 199200 102472
rect 880 96496 199200 96768
rect 880 96488 199120 96496
rect 800 96216 199120 96488
rect 800 90240 199200 96216
rect 800 90104 199120 90240
rect 880 89960 199120 90104
rect 880 89824 199200 89960
rect 800 83984 199200 89824
rect 800 83704 199120 83984
rect 800 83440 199200 83704
rect 880 83160 199200 83440
rect 800 77864 199200 83160
rect 800 77584 199120 77864
rect 800 76776 199200 77584
rect 880 76496 199200 76776
rect 800 71608 199200 76496
rect 800 71328 199120 71608
rect 800 70112 199200 71328
rect 880 69832 199200 70112
rect 800 65352 199200 69832
rect 800 65072 199120 65352
rect 800 63448 199200 65072
rect 880 63168 199200 63448
rect 800 59096 199200 63168
rect 800 58816 199120 59096
rect 800 56784 199200 58816
rect 880 56504 199200 56784
rect 800 52976 199200 56504
rect 800 52696 199120 52976
rect 800 50120 199200 52696
rect 880 49840 199200 50120
rect 800 46720 199200 49840
rect 800 46440 199120 46720
rect 800 43456 199200 46440
rect 880 43176 199200 43456
rect 800 40464 199200 43176
rect 800 40184 199120 40464
rect 800 36792 199200 40184
rect 880 36512 199200 36792
rect 800 34208 199200 36512
rect 800 33928 199120 34208
rect 800 30128 199200 33928
rect 880 29848 199200 30128
rect 800 28088 199200 29848
rect 800 27808 199120 28088
rect 800 23464 199200 27808
rect 880 23184 199200 23464
rect 800 21832 199200 23184
rect 800 21552 199120 21832
rect 800 16800 199200 21552
rect 880 16520 199200 16800
rect 800 15576 199200 16520
rect 800 15296 199120 15576
rect 800 10136 199200 15296
rect 880 9856 199200 10136
rect 800 9320 199200 9856
rect 800 9040 199120 9320
rect 800 3472 199200 9040
rect 880 3200 199200 3472
rect 880 3192 199120 3200
rect 800 2920 199120 3192
rect 800 2143 199200 2920
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
<< obsm4 >>
rect 20483 2347 34848 70549
rect 35328 2347 50208 70549
rect 50688 2347 65568 70549
rect 66048 2347 80928 70549
rect 81408 2347 90653 70549
<< labels >>
rlabel metal3 s 199200 3000 200000 3120 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 199200 189592 200000 189712 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 199200 208224 200000 208344 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 199200 226992 200000 227112 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 199200 245624 200000 245744 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 199200 264256 200000 264376 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 196254 279200 196310 280000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 173990 279200 174046 280000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 151818 279200 151874 280000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 129554 279200 129610 280000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 107382 279200 107438 280000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 199200 21632 200000 21752 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 85118 279200 85174 280000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 62946 279200 63002 280000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 40682 279200 40738 280000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 18510 279200 18566 280000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 276496 800 276616 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 256504 800 256624 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 236512 800 236632 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 216520 800 216640 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 176536 800 176656 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 199200 40264 200000 40384 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 199200 58896 200000 59016 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 199200 77664 200000 77784 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 199200 96296 200000 96416 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 199200 114928 200000 115048 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 199200 133560 200000 133680 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 199200 152328 200000 152448 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 199200 170960 200000 171080 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 199200 15376 200000 15496 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 199200 202104 200000 202224 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 199200 220736 200000 220856 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 199200 239368 200000 239488 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 199200 258000 200000 258120 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 199200 276768 200000 276888 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 181442 279200 181498 280000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 159178 279200 159234 280000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 137006 279200 137062 280000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 114742 279200 114798 280000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92570 279200 92626 280000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 199200 34008 200000 34128 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 70306 279200 70362 280000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 48134 279200 48190 280000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 25870 279200 25926 280000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 3698 279200 3754 280000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 263168 800 263288 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 243176 800 243296 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 223184 800 223304 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 203192 800 203312 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 183200 800 183320 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 163208 800 163328 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 199200 52776 200000 52896 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 143216 800 143336 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 199200 71408 200000 71528 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 199200 90040 200000 90160 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 199200 108672 200000 108792 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 199200 127440 200000 127560 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 199200 146072 200000 146192 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 199200 164704 200000 164824 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 199200 183336 200000 183456 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 199200 9120 200000 9240 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 199200 195848 200000 195968 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 199200 214480 200000 214600 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 199200 233112 200000 233232 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 199200 251880 200000 252000 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 199200 270512 200000 270632 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 188802 279200 188858 280000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 166630 279200 166686 280000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 144366 279200 144422 280000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 122194 279200 122250 280000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 99930 279200 99986 280000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 199200 27888 200000 28008 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 77758 279200 77814 280000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 55494 279200 55550 280000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 33322 279200 33378 280000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 11058 279200 11114 280000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 269832 800 269952 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 249840 800 249960 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 229848 800 229968 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 209856 800 209976 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 189864 800 189984 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 169872 800 169992 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 199200 46520 200000 46640 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 149880 800 150000 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 199200 65152 200000 65272 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 199200 83784 200000 83904 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 199200 102552 200000 102672 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 199200 121184 200000 121304 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 199200 139816 200000 139936 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 199200 158448 200000 158568 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 199200 177216 200000 177336 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 199382 0 199438 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 166446 0 166502 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 181074 0 181130 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 184754 0 184810 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 189630 0 189686 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 192022 0 192078 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 193310 0 193366 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 194506 0 194562 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 164054 0 164110 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26987970
string GDS_FILE /home/tutel/caravel_tutorial/RNG-SCROLL/openlane/user_proj_example/runs/user_proj_example/results/signoff/user_proj_example.magic.gds
string GDS_START 1388334
<< end >>

