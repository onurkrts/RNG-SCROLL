magic
tech sky130A
magscale 1 2
timestamp 1654504549
<< obsli1 >>
rect 1104 2159 158884 237745
<< obsm1 >>
rect 106 960 159790 237776
<< metal2 >>
rect 2962 239200 3018 240000
rect 8850 239200 8906 240000
rect 14738 239200 14794 240000
rect 20718 239200 20774 240000
rect 26606 239200 26662 240000
rect 32586 239200 32642 240000
rect 38474 239200 38530 240000
rect 44362 239200 44418 240000
rect 50342 239200 50398 240000
rect 56230 239200 56286 240000
rect 62210 239200 62266 240000
rect 68098 239200 68154 240000
rect 73986 239200 74042 240000
rect 79966 239200 80022 240000
rect 85854 239200 85910 240000
rect 91834 239200 91890 240000
rect 97722 239200 97778 240000
rect 103610 239200 103666 240000
rect 109590 239200 109646 240000
rect 115478 239200 115534 240000
rect 121458 239200 121514 240000
rect 127346 239200 127402 240000
rect 133234 239200 133290 240000
rect 139214 239200 139270 240000
rect 145102 239200 145158 240000
rect 151082 239200 151138 240000
rect 156970 239200 157026 240000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159362 0 159418 800
rect 159730 0 159786 800
<< obsm2 >>
rect 112 239144 2906 239306
rect 3074 239144 8794 239306
rect 8962 239144 14682 239306
rect 14850 239144 20662 239306
rect 20830 239144 26550 239306
rect 26718 239144 32530 239306
rect 32698 239144 38418 239306
rect 38586 239144 44306 239306
rect 44474 239144 50286 239306
rect 50454 239144 56174 239306
rect 56342 239144 62154 239306
rect 62322 239144 68042 239306
rect 68210 239144 73930 239306
rect 74098 239144 79910 239306
rect 80078 239144 85798 239306
rect 85966 239144 91778 239306
rect 91946 239144 97666 239306
rect 97834 239144 103554 239306
rect 103722 239144 109534 239306
rect 109702 239144 115422 239306
rect 115590 239144 121402 239306
rect 121570 239144 127290 239306
rect 127458 239144 133178 239306
rect 133346 239144 139158 239306
rect 139326 239144 145046 239306
rect 145214 239144 151026 239306
rect 151194 239144 156914 239306
rect 157082 239144 159784 239306
rect 112 856 159784 239144
rect 222 734 330 856
rect 498 734 698 856
rect 866 734 974 856
rect 1142 734 1342 856
rect 1510 734 1618 856
rect 1786 734 1986 856
rect 2154 734 2262 856
rect 2430 734 2630 856
rect 2798 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3550 856
rect 3718 734 3918 856
rect 4086 734 4194 856
rect 4362 734 4562 856
rect 4730 734 4838 856
rect 5006 734 5206 856
rect 5374 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6494 856
rect 6662 734 6862 856
rect 7030 734 7138 856
rect 7306 734 7506 856
rect 7674 734 7782 856
rect 7950 734 8150 856
rect 8318 734 8426 856
rect 8594 734 8794 856
rect 8962 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9714 856
rect 9882 734 10082 856
rect 10250 734 10358 856
rect 10526 734 10726 856
rect 10894 734 11002 856
rect 11170 734 11370 856
rect 11538 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12658 856
rect 12826 734 13026 856
rect 13194 734 13302 856
rect 13470 734 13670 856
rect 13838 734 13946 856
rect 14114 734 14314 856
rect 14482 734 14590 856
rect 14758 734 14958 856
rect 15126 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15878 856
rect 16046 734 16246 856
rect 16414 734 16522 856
rect 16690 734 16890 856
rect 17058 734 17166 856
rect 17334 734 17534 856
rect 17702 734 17902 856
rect 18070 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18822 856
rect 18990 734 19190 856
rect 19358 734 19466 856
rect 19634 734 19834 856
rect 20002 734 20110 856
rect 20278 734 20478 856
rect 20646 734 20754 856
rect 20922 734 21122 856
rect 21290 734 21398 856
rect 21566 734 21766 856
rect 21934 734 22042 856
rect 22210 734 22410 856
rect 22578 734 22686 856
rect 22854 734 23054 856
rect 23222 734 23330 856
rect 23498 734 23698 856
rect 23866 734 24066 856
rect 24234 734 24342 856
rect 24510 734 24710 856
rect 24878 734 24986 856
rect 25154 734 25354 856
rect 25522 734 25630 856
rect 25798 734 25998 856
rect 26166 734 26274 856
rect 26442 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27562 856
rect 27730 734 27930 856
rect 28098 734 28206 856
rect 28374 734 28574 856
rect 28742 734 28850 856
rect 29018 734 29218 856
rect 29386 734 29494 856
rect 29662 734 29862 856
rect 30030 734 30230 856
rect 30398 734 30506 856
rect 30674 734 30874 856
rect 31042 734 31150 856
rect 31318 734 31518 856
rect 31686 734 31794 856
rect 31962 734 32162 856
rect 32330 734 32438 856
rect 32606 734 32806 856
rect 32974 734 33082 856
rect 33250 734 33450 856
rect 33618 734 33726 856
rect 33894 734 34094 856
rect 34262 734 34370 856
rect 34538 734 34738 856
rect 34906 734 35014 856
rect 35182 734 35382 856
rect 35550 734 35750 856
rect 35918 734 36026 856
rect 36194 734 36394 856
rect 36562 734 36670 856
rect 36838 734 37038 856
rect 37206 734 37314 856
rect 37482 734 37682 856
rect 37850 734 37958 856
rect 38126 734 38326 856
rect 38494 734 38602 856
rect 38770 734 38970 856
rect 39138 734 39246 856
rect 39414 734 39614 856
rect 39782 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40534 856
rect 40702 734 40902 856
rect 41070 734 41178 856
rect 41346 734 41546 856
rect 41714 734 41914 856
rect 42082 734 42190 856
rect 42358 734 42558 856
rect 42726 734 42834 856
rect 43002 734 43202 856
rect 43370 734 43478 856
rect 43646 734 43846 856
rect 44014 734 44122 856
rect 44290 734 44490 856
rect 44658 734 44766 856
rect 44934 734 45134 856
rect 45302 734 45410 856
rect 45578 734 45778 856
rect 45946 734 46054 856
rect 46222 734 46422 856
rect 46590 734 46698 856
rect 46866 734 47066 856
rect 47234 734 47342 856
rect 47510 734 47710 856
rect 47878 734 48078 856
rect 48246 734 48354 856
rect 48522 734 48722 856
rect 48890 734 48998 856
rect 49166 734 49366 856
rect 49534 734 49642 856
rect 49810 734 50010 856
rect 50178 734 50286 856
rect 50454 734 50654 856
rect 50822 734 50930 856
rect 51098 734 51298 856
rect 51466 734 51574 856
rect 51742 734 51942 856
rect 52110 734 52218 856
rect 52386 734 52586 856
rect 52754 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53874 856
rect 54042 734 54242 856
rect 54410 734 54518 856
rect 54686 734 54886 856
rect 55054 734 55162 856
rect 55330 734 55530 856
rect 55698 734 55806 856
rect 55974 734 56174 856
rect 56342 734 56450 856
rect 56618 734 56818 856
rect 56986 734 57094 856
rect 57262 734 57462 856
rect 57630 734 57738 856
rect 57906 734 58106 856
rect 58274 734 58382 856
rect 58550 734 58750 856
rect 58918 734 59026 856
rect 59194 734 59394 856
rect 59562 734 59762 856
rect 59930 734 60038 856
rect 60206 734 60406 856
rect 60574 734 60682 856
rect 60850 734 61050 856
rect 61218 734 61326 856
rect 61494 734 61694 856
rect 61862 734 61970 856
rect 62138 734 62338 856
rect 62506 734 62614 856
rect 62782 734 62982 856
rect 63150 734 63258 856
rect 63426 734 63626 856
rect 63794 734 63902 856
rect 64070 734 64270 856
rect 64438 734 64546 856
rect 64714 734 64914 856
rect 65082 734 65282 856
rect 65450 734 65558 856
rect 65726 734 65926 856
rect 66094 734 66202 856
rect 66370 734 66570 856
rect 66738 734 66846 856
rect 67014 734 67214 856
rect 67382 734 67490 856
rect 67658 734 67858 856
rect 68026 734 68134 856
rect 68302 734 68502 856
rect 68670 734 68778 856
rect 68946 734 69146 856
rect 69314 734 69422 856
rect 69590 734 69790 856
rect 69958 734 70066 856
rect 70234 734 70434 856
rect 70602 734 70710 856
rect 70878 734 71078 856
rect 71246 734 71446 856
rect 71614 734 71722 856
rect 71890 734 72090 856
rect 72258 734 72366 856
rect 72534 734 72734 856
rect 72902 734 73010 856
rect 73178 734 73378 856
rect 73546 734 73654 856
rect 73822 734 74022 856
rect 74190 734 74298 856
rect 74466 734 74666 856
rect 74834 734 74942 856
rect 75110 734 75310 856
rect 75478 734 75586 856
rect 75754 734 75954 856
rect 76122 734 76230 856
rect 76398 734 76598 856
rect 76766 734 76874 856
rect 77042 734 77242 856
rect 77410 734 77610 856
rect 77778 734 77886 856
rect 78054 734 78254 856
rect 78422 734 78530 856
rect 78698 734 78898 856
rect 79066 734 79174 856
rect 79342 734 79542 856
rect 79710 734 79818 856
rect 79986 734 80186 856
rect 80354 734 80462 856
rect 80630 734 80830 856
rect 80998 734 81106 856
rect 81274 734 81474 856
rect 81642 734 81750 856
rect 81918 734 82118 856
rect 82286 734 82394 856
rect 82562 734 82762 856
rect 82930 734 83130 856
rect 83298 734 83406 856
rect 83574 734 83774 856
rect 83942 734 84050 856
rect 84218 734 84418 856
rect 84586 734 84694 856
rect 84862 734 85062 856
rect 85230 734 85338 856
rect 85506 734 85706 856
rect 85874 734 85982 856
rect 86150 734 86350 856
rect 86518 734 86626 856
rect 86794 734 86994 856
rect 87162 734 87270 856
rect 87438 734 87638 856
rect 87806 734 87914 856
rect 88082 734 88282 856
rect 88450 734 88558 856
rect 88726 734 88926 856
rect 89094 734 89294 856
rect 89462 734 89570 856
rect 89738 734 89938 856
rect 90106 734 90214 856
rect 90382 734 90582 856
rect 90750 734 90858 856
rect 91026 734 91226 856
rect 91394 734 91502 856
rect 91670 734 91870 856
rect 92038 734 92146 856
rect 92314 734 92514 856
rect 92682 734 92790 856
rect 92958 734 93158 856
rect 93326 734 93434 856
rect 93602 734 93802 856
rect 93970 734 94078 856
rect 94246 734 94446 856
rect 94614 734 94722 856
rect 94890 734 95090 856
rect 95258 734 95458 856
rect 95626 734 95734 856
rect 95902 734 96102 856
rect 96270 734 96378 856
rect 96546 734 96746 856
rect 96914 734 97022 856
rect 97190 734 97390 856
rect 97558 734 97666 856
rect 97834 734 98034 856
rect 98202 734 98310 856
rect 98478 734 98678 856
rect 98846 734 98954 856
rect 99122 734 99322 856
rect 99490 734 99598 856
rect 99766 734 99966 856
rect 100134 734 100242 856
rect 100410 734 100610 856
rect 100778 734 100978 856
rect 101146 734 101254 856
rect 101422 734 101622 856
rect 101790 734 101898 856
rect 102066 734 102266 856
rect 102434 734 102542 856
rect 102710 734 102910 856
rect 103078 734 103186 856
rect 103354 734 103554 856
rect 103722 734 103830 856
rect 103998 734 104198 856
rect 104366 734 104474 856
rect 104642 734 104842 856
rect 105010 734 105118 856
rect 105286 734 105486 856
rect 105654 734 105762 856
rect 105930 734 106130 856
rect 106298 734 106406 856
rect 106574 734 106774 856
rect 106942 734 107142 856
rect 107310 734 107418 856
rect 107586 734 107786 856
rect 107954 734 108062 856
rect 108230 734 108430 856
rect 108598 734 108706 856
rect 108874 734 109074 856
rect 109242 734 109350 856
rect 109518 734 109718 856
rect 109886 734 109994 856
rect 110162 734 110362 856
rect 110530 734 110638 856
rect 110806 734 111006 856
rect 111174 734 111282 856
rect 111450 734 111650 856
rect 111818 734 111926 856
rect 112094 734 112294 856
rect 112462 734 112662 856
rect 112830 734 112938 856
rect 113106 734 113306 856
rect 113474 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114226 856
rect 114394 734 114594 856
rect 114762 734 114870 856
rect 115038 734 115238 856
rect 115406 734 115514 856
rect 115682 734 115882 856
rect 116050 734 116158 856
rect 116326 734 116526 856
rect 116694 734 116802 856
rect 116970 734 117170 856
rect 117338 734 117446 856
rect 117614 734 117814 856
rect 117982 734 118090 856
rect 118258 734 118458 856
rect 118626 734 118826 856
rect 118994 734 119102 856
rect 119270 734 119470 856
rect 119638 734 119746 856
rect 119914 734 120114 856
rect 120282 734 120390 856
rect 120558 734 120758 856
rect 120926 734 121034 856
rect 121202 734 121402 856
rect 121570 734 121678 856
rect 121846 734 122046 856
rect 122214 734 122322 856
rect 122490 734 122690 856
rect 122858 734 122966 856
rect 123134 734 123334 856
rect 123502 734 123610 856
rect 123778 734 123978 856
rect 124146 734 124254 856
rect 124422 734 124622 856
rect 124790 734 124990 856
rect 125158 734 125266 856
rect 125434 734 125634 856
rect 125802 734 125910 856
rect 126078 734 126278 856
rect 126446 734 126554 856
rect 126722 734 126922 856
rect 127090 734 127198 856
rect 127366 734 127566 856
rect 127734 734 127842 856
rect 128010 734 128210 856
rect 128378 734 128486 856
rect 128654 734 128854 856
rect 129022 734 129130 856
rect 129298 734 129498 856
rect 129666 734 129774 856
rect 129942 734 130142 856
rect 130310 734 130510 856
rect 130678 734 130786 856
rect 130954 734 131154 856
rect 131322 734 131430 856
rect 131598 734 131798 856
rect 131966 734 132074 856
rect 132242 734 132442 856
rect 132610 734 132718 856
rect 132886 734 133086 856
rect 133254 734 133362 856
rect 133530 734 133730 856
rect 133898 734 134006 856
rect 134174 734 134374 856
rect 134542 734 134650 856
rect 134818 734 135018 856
rect 135186 734 135294 856
rect 135462 734 135662 856
rect 135830 734 135938 856
rect 136106 734 136306 856
rect 136474 734 136674 856
rect 136842 734 136950 856
rect 137118 734 137318 856
rect 137486 734 137594 856
rect 137762 734 137962 856
rect 138130 734 138238 856
rect 138406 734 138606 856
rect 138774 734 138882 856
rect 139050 734 139250 856
rect 139418 734 139526 856
rect 139694 734 139894 856
rect 140062 734 140170 856
rect 140338 734 140538 856
rect 140706 734 140814 856
rect 140982 734 141182 856
rect 141350 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142102 856
rect 142270 734 142470 856
rect 142638 734 142838 856
rect 143006 734 143114 856
rect 143282 734 143482 856
rect 143650 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144402 856
rect 144570 734 144770 856
rect 144938 734 145046 856
rect 145214 734 145414 856
rect 145582 734 145690 856
rect 145858 734 146058 856
rect 146226 734 146334 856
rect 146502 734 146702 856
rect 146870 734 146978 856
rect 147146 734 147346 856
rect 147514 734 147622 856
rect 147790 734 147990 856
rect 148158 734 148358 856
rect 148526 734 148634 856
rect 148802 734 149002 856
rect 149170 734 149278 856
rect 149446 734 149646 856
rect 149814 734 149922 856
rect 150090 734 150290 856
rect 150458 734 150566 856
rect 150734 734 150934 856
rect 151102 734 151210 856
rect 151378 734 151578 856
rect 151746 734 151854 856
rect 152022 734 152222 856
rect 152390 734 152498 856
rect 152666 734 152866 856
rect 153034 734 153142 856
rect 153310 734 153510 856
rect 153678 734 153786 856
rect 153954 734 154154 856
rect 154322 734 154522 856
rect 154690 734 154798 856
rect 154966 734 155166 856
rect 155334 734 155442 856
rect 155610 734 155810 856
rect 155978 734 156086 856
rect 156254 734 156454 856
rect 156622 734 156730 856
rect 156898 734 157098 856
rect 157266 734 157374 856
rect 157542 734 157742 856
rect 157910 734 158018 856
rect 158186 734 158386 856
rect 158554 734 158662 856
rect 158830 734 159030 856
rect 159198 734 159306 856
rect 159474 734 159674 856
<< metal3 >>
rect 0 237056 800 237176
rect 159200 237192 160000 237312
rect 159200 231888 160000 232008
rect 0 231344 800 231464
rect 159200 226584 160000 226704
rect 0 225632 800 225752
rect 159200 221280 160000 221400
rect 0 219920 800 220040
rect 159200 215840 160000 215960
rect 0 214208 800 214328
rect 159200 210536 160000 210656
rect 0 208496 800 208616
rect 159200 205232 160000 205352
rect 0 202784 800 202904
rect 159200 199928 160000 200048
rect 0 197072 800 197192
rect 159200 194624 160000 194744
rect 0 191360 800 191480
rect 159200 189184 160000 189304
rect 0 185648 800 185768
rect 159200 183880 160000 184000
rect 0 179936 800 180056
rect 159200 178576 160000 178696
rect 0 174224 800 174344
rect 159200 173272 160000 173392
rect 0 168512 800 168632
rect 159200 167832 160000 167952
rect 0 162800 800 162920
rect 159200 162528 160000 162648
rect 0 157088 800 157208
rect 159200 157224 160000 157344
rect 159200 151920 160000 152040
rect 0 151376 800 151496
rect 159200 146616 160000 146736
rect 0 145664 800 145784
rect 159200 141176 160000 141296
rect 0 139952 800 140072
rect 159200 135872 160000 135992
rect 0 134240 800 134360
rect 159200 130568 160000 130688
rect 0 128528 800 128648
rect 159200 125264 160000 125384
rect 0 122816 800 122936
rect 159200 119824 160000 119944
rect 0 117104 800 117224
rect 159200 114520 160000 114640
rect 0 111392 800 111512
rect 159200 109216 160000 109336
rect 0 105680 800 105800
rect 159200 103912 160000 104032
rect 0 99968 800 100088
rect 159200 98608 160000 98728
rect 0 94256 800 94376
rect 159200 93168 160000 93288
rect 0 88544 800 88664
rect 159200 87864 160000 87984
rect 0 82832 800 82952
rect 159200 82560 160000 82680
rect 0 77120 800 77240
rect 159200 77256 160000 77376
rect 159200 71816 160000 71936
rect 0 71408 800 71528
rect 159200 66512 160000 66632
rect 0 65696 800 65816
rect 159200 61208 160000 61328
rect 0 59984 800 60104
rect 159200 55904 160000 56024
rect 0 54272 800 54392
rect 159200 50600 160000 50720
rect 0 48560 800 48680
rect 159200 45160 160000 45280
rect 0 42848 800 42968
rect 159200 39856 160000 39976
rect 0 37136 800 37256
rect 159200 34552 160000 34672
rect 0 31424 800 31544
rect 159200 29248 160000 29368
rect 0 25712 800 25832
rect 159200 23808 160000 23928
rect 0 20000 800 20120
rect 159200 18504 160000 18624
rect 0 14288 800 14408
rect 159200 13200 160000 13320
rect 0 8576 800 8696
rect 159200 7896 160000 8016
rect 0 2864 800 2984
rect 159200 2592 160000 2712
<< obsm3 >>
rect 800 237392 159200 237761
rect 800 237256 159120 237392
rect 880 237112 159120 237256
rect 880 236976 159200 237112
rect 800 232088 159200 236976
rect 800 231808 159120 232088
rect 800 231544 159200 231808
rect 880 231264 159200 231544
rect 800 226784 159200 231264
rect 800 226504 159120 226784
rect 800 225832 159200 226504
rect 880 225552 159200 225832
rect 800 221480 159200 225552
rect 800 221200 159120 221480
rect 800 220120 159200 221200
rect 880 219840 159200 220120
rect 800 216040 159200 219840
rect 800 215760 159120 216040
rect 800 214408 159200 215760
rect 880 214128 159200 214408
rect 800 210736 159200 214128
rect 800 210456 159120 210736
rect 800 208696 159200 210456
rect 880 208416 159200 208696
rect 800 205432 159200 208416
rect 800 205152 159120 205432
rect 800 202984 159200 205152
rect 880 202704 159200 202984
rect 800 200128 159200 202704
rect 800 199848 159120 200128
rect 800 197272 159200 199848
rect 880 196992 159200 197272
rect 800 194824 159200 196992
rect 800 194544 159120 194824
rect 800 191560 159200 194544
rect 880 191280 159200 191560
rect 800 189384 159200 191280
rect 800 189104 159120 189384
rect 800 185848 159200 189104
rect 880 185568 159200 185848
rect 800 184080 159200 185568
rect 800 183800 159120 184080
rect 800 180136 159200 183800
rect 880 179856 159200 180136
rect 800 178776 159200 179856
rect 800 178496 159120 178776
rect 800 174424 159200 178496
rect 880 174144 159200 174424
rect 800 173472 159200 174144
rect 800 173192 159120 173472
rect 800 168712 159200 173192
rect 880 168432 159200 168712
rect 800 168032 159200 168432
rect 800 167752 159120 168032
rect 800 163000 159200 167752
rect 880 162728 159200 163000
rect 880 162720 159120 162728
rect 800 162448 159120 162720
rect 800 157424 159200 162448
rect 800 157288 159120 157424
rect 880 157144 159120 157288
rect 880 157008 159200 157144
rect 800 152120 159200 157008
rect 800 151840 159120 152120
rect 800 151576 159200 151840
rect 880 151296 159200 151576
rect 800 146816 159200 151296
rect 800 146536 159120 146816
rect 800 145864 159200 146536
rect 880 145584 159200 145864
rect 800 141376 159200 145584
rect 800 141096 159120 141376
rect 800 140152 159200 141096
rect 880 139872 159200 140152
rect 800 136072 159200 139872
rect 800 135792 159120 136072
rect 800 134440 159200 135792
rect 880 134160 159200 134440
rect 800 130768 159200 134160
rect 800 130488 159120 130768
rect 800 128728 159200 130488
rect 880 128448 159200 128728
rect 800 125464 159200 128448
rect 800 125184 159120 125464
rect 800 123016 159200 125184
rect 880 122736 159200 123016
rect 800 120024 159200 122736
rect 800 119744 159120 120024
rect 800 117304 159200 119744
rect 880 117024 159200 117304
rect 800 114720 159200 117024
rect 800 114440 159120 114720
rect 800 111592 159200 114440
rect 880 111312 159200 111592
rect 800 109416 159200 111312
rect 800 109136 159120 109416
rect 800 105880 159200 109136
rect 880 105600 159200 105880
rect 800 104112 159200 105600
rect 800 103832 159120 104112
rect 800 100168 159200 103832
rect 880 99888 159200 100168
rect 800 98808 159200 99888
rect 800 98528 159120 98808
rect 800 94456 159200 98528
rect 880 94176 159200 94456
rect 800 93368 159200 94176
rect 800 93088 159120 93368
rect 800 88744 159200 93088
rect 880 88464 159200 88744
rect 800 88064 159200 88464
rect 800 87784 159120 88064
rect 800 83032 159200 87784
rect 880 82760 159200 83032
rect 880 82752 159120 82760
rect 800 82480 159120 82752
rect 800 77456 159200 82480
rect 800 77320 159120 77456
rect 880 77176 159120 77320
rect 880 77040 159200 77176
rect 800 72016 159200 77040
rect 800 71736 159120 72016
rect 800 71608 159200 71736
rect 880 71328 159200 71608
rect 800 66712 159200 71328
rect 800 66432 159120 66712
rect 800 65896 159200 66432
rect 880 65616 159200 65896
rect 800 61408 159200 65616
rect 800 61128 159120 61408
rect 800 60184 159200 61128
rect 880 59904 159200 60184
rect 800 56104 159200 59904
rect 800 55824 159120 56104
rect 800 54472 159200 55824
rect 880 54192 159200 54472
rect 800 50800 159200 54192
rect 800 50520 159120 50800
rect 800 48760 159200 50520
rect 880 48480 159200 48760
rect 800 45360 159200 48480
rect 800 45080 159120 45360
rect 800 43048 159200 45080
rect 880 42768 159200 43048
rect 800 40056 159200 42768
rect 800 39776 159120 40056
rect 800 37336 159200 39776
rect 880 37056 159200 37336
rect 800 34752 159200 37056
rect 800 34472 159120 34752
rect 800 31624 159200 34472
rect 880 31344 159200 31624
rect 800 29448 159200 31344
rect 800 29168 159120 29448
rect 800 25912 159200 29168
rect 880 25632 159200 25912
rect 800 24008 159200 25632
rect 800 23728 159120 24008
rect 800 20200 159200 23728
rect 880 19920 159200 20200
rect 800 18704 159200 19920
rect 800 18424 159120 18704
rect 800 14488 159200 18424
rect 880 14208 159200 14488
rect 800 13400 159200 14208
rect 800 13120 159120 13400
rect 800 8776 159200 13120
rect 880 8496 159200 8776
rect 800 8096 159200 8496
rect 800 7816 159120 8096
rect 800 3064 159200 7816
rect 880 2792 159200 3064
rect 880 2784 159120 2792
rect 800 2512 159120 2784
rect 800 2143 159200 2512
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
rect 81008 2128 81328 237776
rect 96368 2128 96688 237776
rect 111728 2128 112048 237776
rect 127088 2128 127408 237776
rect 142448 2128 142768 237776
rect 157808 2128 158128 237776
<< obsm4 >>
rect 19379 2755 19488 89861
rect 19968 2755 34848 89861
rect 35328 2755 50208 89861
rect 50688 2755 65568 89861
rect 66048 2755 76117 89861
<< labels >>
rlabel metal3 s 159200 2592 160000 2712 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 159200 162528 160000 162648 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 159200 178576 160000 178696 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 159200 194624 160000 194744 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 159200 210536 160000 210656 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 159200 226584 160000 226704 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 156970 239200 157026 240000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 139214 239200 139270 240000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 121458 239200 121514 240000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 103610 239200 103666 240000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 85854 239200 85910 240000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 159200 18504 160000 18624 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 68098 239200 68154 240000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50342 239200 50398 240000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 32586 239200 32642 240000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 14738 239200 14794 240000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 237056 800 237176 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 219920 800 220040 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 202784 800 202904 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 151376 800 151496 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 159200 34552 160000 34672 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 159200 50600 160000 50720 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 159200 66512 160000 66632 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 159200 82560 160000 82680 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 159200 98608 160000 98728 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 159200 114520 160000 114640 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 159200 130568 160000 130688 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 159200 146616 160000 146736 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 159200 13200 160000 13320 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 159200 173272 160000 173392 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 159200 189184 160000 189304 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 159200 205232 160000 205352 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 159200 221280 160000 221400 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 159200 237192 160000 237312 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 145102 239200 145158 240000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 127346 239200 127402 240000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 109590 239200 109646 240000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 91834 239200 91890 240000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 73986 239200 74042 240000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 159200 29248 160000 29368 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 56230 239200 56286 240000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 38474 239200 38530 240000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 20718 239200 20774 240000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 2962 239200 3018 240000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 225632 800 225752 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 208496 800 208616 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 191360 800 191480 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 174224 800 174344 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 139952 800 140072 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 159200 45160 160000 45280 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 105680 800 105800 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 159200 61208 160000 61328 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 159200 77256 160000 77376 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 159200 93168 160000 93288 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 159200 109216 160000 109336 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 159200 125264 160000 125384 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 159200 141176 160000 141296 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 159200 157224 160000 157344 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 159200 7896 160000 8016 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 159200 167832 160000 167952 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 159200 183880 160000 184000 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 159200 199928 160000 200048 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 159200 215840 160000 215960 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 159200 231888 160000 232008 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 151082 239200 151138 240000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 133234 239200 133290 240000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 115478 239200 115534 240000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 97722 239200 97778 240000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 79966 239200 80022 240000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 159200 23808 160000 23928 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 62210 239200 62266 240000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 44362 239200 44418 240000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 26606 239200 26662 240000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 8850 239200 8906 240000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 231344 800 231464 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 179936 800 180056 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 162800 800 162920 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 145664 800 145784 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 159200 39856 160000 39976 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 159200 55904 160000 56024 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 159200 71816 160000 71936 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 159200 87864 160000 87984 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 159200 103912 160000 104032 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 159200 119824 160000 119944 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 159200 135872 160000 135992 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 159200 151920 160000 152040 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 159730 0 159786 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 160000 240000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22324538
string GDS_FILE /home/tutel/caravel_tutorial/RNG-SCROLL/openlane/user_proj_example/runs/user_proj_example/results/signoff/user_proj_example.magic.gds
string GDS_START 1284618
<< end >>

